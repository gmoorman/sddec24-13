magic
tech sky130B
magscale 1 2
timestamp 1733718626
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 183
rect 29 -17 63 21
<< scnmos >>
rect 79 47 657 157
<< scpmoshvt >>
rect 79 323 657 497
<< ndiff >>
rect 27 112 79 157
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 657 112 709 157
rect 657 78 667 112
rect 701 78 709 112
rect 657 47 709 78
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 383 79 451
rect 27 349 35 383
rect 69 349 79 383
rect 27 323 79 349
rect 657 485 709 497
rect 657 451 667 485
rect 701 451 709 485
rect 657 383 709 451
rect 657 349 667 383
rect 701 349 709 383
rect 657 323 709 349
<< ndiffc >>
rect 35 78 69 112
rect 667 78 701 112
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 667 451 701 485
rect 667 349 701 383
<< poly >>
rect 79 497 657 523
rect 79 297 657 323
rect 79 275 343 297
rect 79 241 95 275
rect 129 241 194 275
rect 228 241 293 275
rect 327 241 343 275
rect 79 225 343 241
rect 385 239 657 255
rect 385 205 401 239
rect 435 205 504 239
rect 538 205 607 239
rect 641 205 657 239
rect 385 183 657 205
rect 79 157 657 183
rect 79 21 657 47
<< polycont >>
rect 95 241 129 275
rect 194 241 228 275
rect 293 241 327 275
rect 401 205 435 239
rect 504 205 538 239
rect 607 205 641 239
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 485 719 527
rect 17 451 35 485
rect 69 451 667 485
rect 701 451 719 485
rect 17 383 719 451
rect 17 349 35 383
rect 69 349 667 383
rect 701 349 719 383
rect 17 309 719 349
rect 17 241 95 275
rect 129 241 194 275
rect 228 241 293 275
rect 327 241 347 275
rect 17 171 347 241
rect 381 239 719 309
rect 381 205 401 239
rect 435 205 504 239
rect 538 205 607 239
rect 641 205 719 239
rect 17 112 719 171
rect 17 78 35 112
rect 69 78 667 112
rect 701 78 719 112
rect 17 17 719 78
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 decap_8
<< properties >>
string FIXED_BBOX 0 0 736 544
string path 0.000 0.000 3.680 0.000 
<< end >>
