magic
tech sky130B
magscale 1 2
timestamp 1731865869
<< metal1 >>
rect 1382 -4362 1418 -4028
rect 1458 -4118 1510 -4108
rect 1458 -4180 1510 -4170
rect 1458 -4450 1494 -4180
rect 1578 -4210 1630 -4200
rect 1578 -4272 1630 -4262
rect 1460 -4492 1494 -4450
rect 1584 -4494 1620 -4272
rect 1662 -4362 1698 -4028
rect 1820 -4118 1872 -4108
rect 1820 -4180 1872 -4170
rect 1304 -5028 1340 -4758
rect 1382 -4924 1418 -4838
rect 1480 -4872 1698 -4838
rect 1374 -4934 1426 -4924
rect 1374 -4996 1426 -4986
rect 1296 -5038 1348 -5028
rect 1480 -5032 1514 -4872
rect 1654 -4934 1706 -4924
rect 1654 -4996 1706 -4986
rect 1296 -5100 1348 -5090
rect 1382 -5066 1514 -5032
rect 1382 -5184 1418 -5066
rect 1458 -5118 1510 -5108
rect 1458 -5180 1510 -5170
rect 1458 -5296 1494 -5180
rect 1662 -5182 1698 -4996
rect 1740 -5014 1776 -4754
rect 1734 -5024 1786 -5014
rect 1734 -5086 1786 -5076
rect 1338 -5814 1374 -5642
rect 1584 -5718 1620 -5482
rect 1706 -5694 1742 -5482
rect 1822 -5694 1872 -4180
rect 1576 -5728 1628 -5718
rect 1706 -5730 1872 -5694
rect 1576 -5790 1628 -5780
rect 1330 -5824 1382 -5814
rect 1330 -5886 1382 -5876
rect 1338 -6014 1374 -5886
rect 1584 -6014 1620 -5790
<< via1 >>
rect 1458 -4170 1510 -4118
rect 1578 -4262 1630 -4210
rect 1820 -4170 1872 -4118
rect 1374 -4986 1426 -4934
rect 1654 -4986 1706 -4934
rect 1296 -5090 1348 -5038
rect 1458 -5170 1510 -5118
rect 1734 -5076 1786 -5024
rect 1576 -5780 1628 -5728
rect 1330 -5876 1382 -5824
<< metal2 >>
rect 1448 -4170 1458 -4118
rect 1510 -4170 1820 -4118
rect 1872 -4170 1882 -4118
rect 1568 -4262 1578 -4210
rect 1630 -4262 1876 -4210
rect 1364 -4986 1374 -4934
rect 1426 -4986 1654 -4934
rect 1706 -4986 1716 -4934
rect 1724 -5036 1734 -5024
rect 1286 -5090 1296 -5038
rect 1348 -5090 1358 -5038
rect 1554 -5070 1734 -5036
rect 1296 -5728 1348 -5090
rect 1554 -5118 1588 -5070
rect 1724 -5076 1734 -5070
rect 1786 -5076 1796 -5024
rect 1448 -5170 1458 -5118
rect 1510 -5170 1588 -5118
rect 1296 -5780 1576 -5728
rect 1628 -5780 1638 -5728
rect 1826 -5824 1876 -4262
rect 1320 -5876 1330 -5824
rect 1382 -5876 1876 -5824
use sky130_fd_pr__nfet_01v8_PHZV97  xm45
timestamp 1731864020
transform 1 0 1400 0 1 -4600
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm46
timestamp 1731864020
transform 1 0 1680 0 1 -4600
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_72KZQ8  xm47
timestamp 1731864020
transform 1 0 1399 0 1 -5427
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm48
timestamp 1731864020
transform 1 0 1679 0 1 -5427
box -73 -257 73 257
<< end >>
