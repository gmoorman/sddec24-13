* NGSPICE file created from 1T1R.ext - technology: sky130B

.subckt x1T1R SL VSS WL BL
X0 BL XR1.BE sky130_fd_pr_reram__reram_cell area_ox=1
X1 XR1.BE WL.t0 SL.t0 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=0.5
R0 WL WL.t0 273.483
R1 SL SL.t0 23.767
R2 VSS.n5 VSS.n3 3546.67
R3 VSS.n8 VSS.n2 3546.67
R4 VSS.n7 VSS.n3 356.945
R5 VSS.n6 VSS.n2 356.945
R6 VSS.n4 VSS.n0 229.12
R7 VSS.n4 VSS.n1 228.268
R8 VSS.n9 VSS.n1 194.666
R9 VSS.n10 VSS.n0 190.249
R10 VSS.n5 VSS.n4 146.25
R11 VSS.n9 VSS.n8 146.25
R12 VSS.n8 VSS.n7 126.323
R13 VSS.n6 VSS.n5 126.323
R14 VSS.n2 VSS.n0 24.3755
R15 VSS.n3 VSS.n1 24.3755
R16 VSS.n7 VSS.t0 14.7199
R17 VSS.t0 VSS.n6 14.7199
R18 VSS.n10 VSS.n9 4.56658
R19 VSS VSS.n10 1.6755
C0 BL WL 0.01281f
C1 XR1.BE WL 0.768937f
C2 BL SL 0.005996f
C3 SL XR1.BE 0.244458f
C4 SL WL 0.786849f
C5 BL XR1.BE 0.116741f
C6 BL VSS 0.439533f
C7 SL VSS 1.40149f
C8 WL VSS 0.774332f
C9 XR1.BE VSS 0.979062f
.ends

