magic
tech sky130B
magscale 1 2
timestamp 1733216309
<< error_p >>
rect -29 -207 29 -201
rect -29 -241 -17 -207
rect -29 -247 29 -241
<< pwell >>
rect -99 -195 99 257
<< nmos >>
rect -15 -169 15 231
<< ndiff >>
rect -73 218 -15 231
rect -73 184 -61 218
rect -27 184 -15 218
rect -73 150 -15 184
rect -73 116 -61 150
rect -27 116 -15 150
rect -73 82 -15 116
rect -73 48 -61 82
rect -27 48 -15 82
rect -73 14 -15 48
rect -73 -20 -61 14
rect -27 -20 -15 14
rect -73 -54 -15 -20
rect -73 -88 -61 -54
rect -27 -88 -15 -54
rect -73 -122 -15 -88
rect -73 -156 -61 -122
rect -27 -156 -15 -122
rect -73 -169 -15 -156
rect 15 218 73 231
rect 15 184 27 218
rect 61 184 73 218
rect 15 150 73 184
rect 15 116 27 150
rect 61 116 73 150
rect 15 82 73 116
rect 15 48 27 82
rect 61 48 73 82
rect 15 14 73 48
rect 15 -20 27 14
rect 61 -20 73 14
rect 15 -54 73 -20
rect 15 -88 27 -54
rect 61 -88 73 -54
rect 15 -122 73 -88
rect 15 -156 27 -122
rect 61 -156 73 -122
rect 15 -169 73 -156
<< ndiffc >>
rect -61 184 -27 218
rect -61 116 -27 150
rect -61 48 -27 82
rect -61 -20 -27 14
rect -61 -88 -27 -54
rect -61 -156 -27 -122
rect 27 184 61 218
rect 27 116 61 150
rect 27 48 61 82
rect 27 -20 61 14
rect 27 -88 61 -54
rect 27 -156 61 -122
<< poly >>
rect -15 231 15 257
rect -15 -191 15 -169
rect -33 -207 33 -191
rect -33 -241 -17 -207
rect 17 -241 33 -207
rect -33 -257 33 -241
<< polycont >>
rect -17 -241 17 -207
<< locali >>
rect -61 218 -27 235
rect -61 150 -27 158
rect -61 82 -27 86
rect -61 -24 -27 -20
rect -61 -96 -27 -88
rect -61 -173 -27 -156
rect 27 218 61 235
rect 27 150 61 158
rect 27 82 61 86
rect 27 -24 61 -20
rect 27 -96 61 -88
rect 27 -173 61 -156
rect -33 -241 -17 -207
rect 17 -241 33 -207
<< viali >>
rect -61 184 -27 192
rect -61 158 -27 184
rect -61 116 -27 120
rect -61 86 -27 116
rect -61 14 -27 48
rect -61 -54 -27 -24
rect -61 -58 -27 -54
rect -61 -122 -27 -96
rect -61 -130 -27 -122
rect 27 184 61 192
rect 27 158 61 184
rect 27 116 61 120
rect 27 86 61 116
rect 27 14 61 48
rect 27 -54 61 -24
rect 27 -58 61 -54
rect 27 -122 61 -96
rect 27 -130 61 -122
rect -17 -241 17 -207
<< metal1 >>
rect -67 192 -21 231
rect -67 158 -61 192
rect -27 158 -21 192
rect -67 120 -21 158
rect -67 86 -61 120
rect -27 86 -21 120
rect -67 48 -21 86
rect -67 14 -61 48
rect -27 14 -21 48
rect -67 -24 -21 14
rect -67 -58 -61 -24
rect -27 -58 -21 -24
rect -67 -96 -21 -58
rect -67 -130 -61 -96
rect -27 -130 -21 -96
rect -67 -169 -21 -130
rect 21 192 67 231
rect 21 158 27 192
rect 61 158 67 192
rect 21 120 67 158
rect 21 86 27 120
rect 61 86 67 120
rect 21 48 67 86
rect 21 14 27 48
rect 61 14 67 48
rect 21 -24 67 14
rect 21 -58 27 -24
rect 61 -58 67 -24
rect 21 -96 67 -58
rect 21 -130 27 -96
rect 61 -130 67 -96
rect 21 -169 67 -130
rect -29 -207 29 -201
rect -29 -241 -17 -207
rect 17 -241 29 -207
rect -29 -247 29 -241
<< end >>
