magic
tech sky130B
magscale 1 2
timestamp 1733717322
<< xpolycontact >>
rect -50 50 50 482
rect -50 -482 50 -50
<< ppolyres >>
rect -50 -50 50 50
<< viali >>
rect -34 67 34 464
rect -34 -464 34 -67
<< metal1 >>
rect -40 464 40 476
rect -40 67 -34 464
rect 34 67 40 464
rect -40 55 40 67
rect -40 -67 40 -55
rect -40 -464 -34 -67
rect 34 -464 40 -67
rect -40 -476 40 -464
<< properties >>
string gencell sky130_fd_pr__res_high_po_5p73
string library sky130
string parameters w 0.5 l 0.5 m 1 nx 1 wmin 5.730 lmin 0.50 rho 319.8 val 95.905 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 1 full_metal 0 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
