magic
tech sky130B
magscale 1 2
timestamp 1733649010
<< viali >>
rect 3341 5321 3375 5355
rect 5457 5253 5491 5287
rect 2789 5185 2823 5219
rect 2881 5185 2915 5219
rect 3157 5185 3191 5219
rect 3433 5185 3467 5219
rect 3893 5185 3927 5219
rect 4353 5185 4387 5219
rect 4537 5185 4571 5219
rect 4629 5185 4663 5219
rect 4997 5185 5031 5219
rect 5181 5185 5215 5219
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 1593 5117 1627 5151
rect 4813 5117 4847 5151
rect 5089 5117 5123 5151
rect 5274 5117 5308 5151
rect 5549 5117 5583 5151
rect 6101 5117 6135 5151
rect 4077 5049 4111 5083
rect 4445 5049 4479 5083
rect 5917 5049 5951 5083
rect 3065 4981 3099 5015
rect 3617 4981 3651 5015
rect 4169 4981 4203 5015
rect 5457 4981 5491 5015
rect 3617 4777 3651 4811
rect 5273 4777 5307 4811
rect 6285 4709 6319 4743
rect 2145 4641 2179 4675
rect 2697 4573 2731 4607
rect 2881 4573 2915 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 4353 4573 4387 4607
rect 4445 4573 4479 4607
rect 4813 4573 4847 4607
rect 5181 4573 5215 4607
rect 5457 4573 5491 4607
rect 5733 4573 5767 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 6285 4573 6319 4607
rect 6469 4573 6503 4607
rect 4077 4505 4111 4539
rect 4971 4505 5005 4539
rect 3065 4437 3099 4471
rect 3341 4437 3375 4471
rect 5549 4437 5583 4471
rect 4445 4233 4479 4267
rect 5917 4233 5951 4267
rect 3709 4097 3743 4131
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 4905 4097 4939 4131
rect 5089 4097 5123 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 5733 4097 5767 4131
rect 6009 4097 6043 4131
rect 6193 4097 6227 4131
rect 4261 4029 4295 4063
rect 3893 3961 3927 3995
rect 6009 3961 6043 3995
rect 3985 3893 4019 3927
rect 4261 3893 4295 3927
rect 4629 3689 4663 3723
rect 5917 3689 5951 3723
rect 6009 3689 6043 3723
rect 6469 3689 6503 3723
rect 6101 3553 6135 3587
rect 2789 3485 2823 3519
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 4353 3485 4387 3519
rect 4813 3485 4847 3519
rect 4905 3485 4939 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5273 3485 5307 3519
rect 5457 3485 5491 3519
rect 5733 3485 5767 3519
rect 6285 3485 6319 3519
rect 1593 3417 1627 3451
rect 6009 3417 6043 3451
rect 3985 3349 4019 3383
rect 4261 3349 4295 3383
rect 4537 3349 4571 3383
rect 4813 3145 4847 3179
rect 5457 3145 5491 3179
rect 4261 3009 4295 3043
rect 4537 3009 4571 3043
rect 4997 3009 5031 3043
rect 5089 3009 5123 3043
rect 5181 3009 5215 3043
rect 5365 3009 5399 3043
rect 5641 3009 5675 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 4629 2941 4663 2975
rect 4445 2873 4479 2907
rect 5365 2873 5399 2907
rect 4905 2601 4939 2635
rect 6009 2601 6043 2635
rect 4997 2533 5031 2567
rect 5641 2533 5675 2567
rect 2697 2397 2731 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 5273 2397 5307 2431
rect 5457 2397 5491 2431
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 1593 2329 1627 2363
rect 5365 2329 5399 2363
<< metal1 >>
rect 4982 5720 4988 5772
rect 5040 5760 5046 5772
rect 6270 5760 6276 5772
rect 5040 5732 6276 5760
rect 5040 5720 5046 5732
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 3568 5596 5764 5624
rect 3568 5584 3574 5596
rect 5736 5568 5764 5596
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5626 5556 5632 5568
rect 4856 5528 5632 5556
rect 4856 5516 4862 5528
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 1104 5466 6968 5488
rect 1104 5414 2376 5466
rect 2428 5414 2440 5466
rect 2492 5414 2504 5466
rect 2556 5414 2568 5466
rect 2620 5414 2632 5466
rect 2684 5414 3802 5466
rect 3854 5414 3866 5466
rect 3918 5414 3930 5466
rect 3982 5414 3994 5466
rect 4046 5414 4058 5466
rect 4110 5414 5228 5466
rect 5280 5414 5292 5466
rect 5344 5414 5356 5466
rect 5408 5414 5420 5466
rect 5472 5414 5484 5466
rect 5536 5414 6654 5466
rect 6706 5414 6718 5466
rect 6770 5414 6782 5466
rect 6834 5414 6846 5466
rect 6898 5414 6910 5466
rect 6962 5414 6968 5466
rect 1104 5392 6968 5414
rect 3050 5312 3056 5364
rect 3108 5312 3114 5364
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5321 3387 5355
rect 3329 5315 3387 5321
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 3068 5216 3096 5312
rect 2915 5188 3096 5216
rect 3145 5219 3203 5225
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3252 5216 3280 5312
rect 3344 5228 3372 5315
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 6362 5352 6368 5364
rect 3476 5324 6368 5352
rect 3476 5312 3482 5324
rect 3510 5244 3516 5296
rect 3568 5244 3574 5296
rect 3191 5188 3280 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 992 5120 1593 5148
rect 992 5108 998 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 2792 5148 2820 5179
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 3528 5216 3556 5244
rect 3467 5188 3556 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 3878 5176 3884 5228
rect 3936 5176 3942 5228
rect 4356 5225 4384 5324
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 4706 5244 4712 5296
rect 4764 5284 4770 5296
rect 5445 5287 5503 5293
rect 5445 5284 5457 5287
rect 4764 5256 5457 5284
rect 4764 5244 4770 5256
rect 5445 5253 5457 5256
rect 5491 5253 5503 5287
rect 5445 5247 5503 5253
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6454 5284 6460 5296
rect 5592 5256 6460 5284
rect 5592 5244 5598 5256
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4488 5188 4537 5216
rect 4488 5176 4494 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 4890 5216 4896 5228
rect 4663 5188 4896 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 4982 5176 4988 5228
rect 5040 5176 5046 5228
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5736 5225 5764 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 5721 5219 5779 5225
rect 5224 5188 5672 5216
rect 5224 5176 5230 5188
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 2792 5120 4813 5148
rect 1581 5111 1639 5117
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 5074 5108 5080 5160
rect 5132 5108 5138 5160
rect 5262 5151 5320 5157
rect 5262 5117 5274 5151
rect 5308 5117 5320 5151
rect 5262 5111 5320 5117
rect 4065 5083 4123 5089
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 4433 5083 4491 5089
rect 4433 5080 4445 5083
rect 4111 5052 4445 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 4433 5049 4445 5052
rect 4479 5080 4491 5083
rect 4706 5080 4712 5092
rect 4479 5052 4712 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5276 5080 5304 5111
rect 5534 5108 5540 5160
rect 5592 5108 5598 5160
rect 5644 5148 5672 5188
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5994 5176 6000 5228
rect 6052 5176 6058 5228
rect 6181 5220 6239 5225
rect 6181 5219 6408 5220
rect 6181 5185 6193 5219
rect 6227 5216 6408 5219
rect 6546 5216 6552 5228
rect 6227 5192 6552 5216
rect 6227 5185 6239 5192
rect 6380 5188 6552 5192
rect 6181 5179 6239 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5644 5120 6101 5148
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 6089 5111 6147 5117
rect 5350 5080 5356 5092
rect 5276 5052 5356 5080
rect 5350 5040 5356 5052
rect 5408 5080 5414 5092
rect 5905 5083 5963 5089
rect 5905 5080 5917 5083
rect 5408 5052 5917 5080
rect 5408 5040 5414 5052
rect 5905 5049 5917 5052
rect 5951 5049 5963 5083
rect 5905 5043 5963 5049
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 3510 5012 3516 5024
rect 3099 4984 3516 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3602 4972 3608 5024
rect 3660 4972 3666 5024
rect 4154 4972 4160 5024
rect 4212 4972 4218 5024
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 5258 5012 5264 5024
rect 4304 4984 5264 5012
rect 4304 4972 4310 4984
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 5442 4972 5448 5024
rect 5500 4972 5506 5024
rect 1104 4922 6808 4944
rect 1104 4870 1663 4922
rect 1715 4870 1727 4922
rect 1779 4870 1791 4922
rect 1843 4870 1855 4922
rect 1907 4870 1919 4922
rect 1971 4870 3089 4922
rect 3141 4870 3153 4922
rect 3205 4870 3217 4922
rect 3269 4870 3281 4922
rect 3333 4870 3345 4922
rect 3397 4870 4515 4922
rect 4567 4870 4579 4922
rect 4631 4870 4643 4922
rect 4695 4870 4707 4922
rect 4759 4870 4771 4922
rect 4823 4870 5941 4922
rect 5993 4870 6005 4922
rect 6057 4870 6069 4922
rect 6121 4870 6133 4922
rect 6185 4870 6197 4922
rect 6249 4870 6808 4922
rect 1104 4848 6808 4870
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3786 4808 3792 4820
rect 3651 4780 3792 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3786 4768 3792 4780
rect 3844 4808 3850 4820
rect 3844 4780 4384 4808
rect 3844 4768 3850 4780
rect 4356 4752 4384 4780
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 5500 4780 6408 4808
rect 5500 4768 5506 4780
rect 2774 4740 2780 4752
rect 2516 4712 2780 4740
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2516 4672 2544 4712
rect 2774 4700 2780 4712
rect 2832 4700 2838 4752
rect 3326 4700 3332 4752
rect 3384 4740 3390 4752
rect 4062 4740 4068 4752
rect 3384 4712 4068 4740
rect 3384 4700 3390 4712
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 4338 4700 4344 4752
rect 4396 4700 4402 4752
rect 4908 4740 4936 4768
rect 6273 4743 6331 4749
rect 6273 4740 6285 4743
rect 4908 4712 6285 4740
rect 6273 4709 6285 4712
rect 6319 4709 6331 4743
rect 6273 4703 6331 4709
rect 5258 4672 5264 4684
rect 2179 4644 2544 4672
rect 2700 4644 4568 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2700 4613 2728 4644
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 2958 4604 2964 4616
rect 2915 4576 2964 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 3326 4604 3332 4616
rect 3191 4576 3332 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3694 4604 3700 4616
rect 3467 4576 3700 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 4065 4539 4123 4545
rect 4065 4536 4077 4539
rect 2832 4508 4077 4536
rect 2832 4496 2838 4508
rect 4065 4505 4077 4508
rect 4111 4505 4123 4539
rect 4065 4499 4123 4505
rect 3050 4428 3056 4480
rect 3108 4428 3114 4480
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 3418 4468 3424 4480
rect 3375 4440 3424 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 4448 4468 4476 4567
rect 4540 4536 4568 4644
rect 5000 4644 5264 4672
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 5000 4604 5028 4644
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 6380 4672 6408 4780
rect 6288 4644 6408 4672
rect 4856 4576 5028 4604
rect 5169 4607 5227 4613
rect 4856 4564 4862 4576
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5626 4604 5632 4616
rect 5491 4576 5632 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 4959 4539 5017 4545
rect 4959 4536 4971 4539
rect 4540 4508 4971 4536
rect 4959 4505 4971 4508
rect 5005 4505 5017 4539
rect 5177 4536 5205 4567
rect 5626 4564 5632 4576
rect 5684 4604 5690 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5684 4576 5733 4604
rect 5684 4564 5690 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6288 4613 6316 4644
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6196 4536 6224 4567
rect 6362 4564 6368 4616
rect 6420 4564 6426 4616
rect 6454 4564 6460 4616
rect 6512 4564 6518 4616
rect 6380 4536 6408 4564
rect 5177 4508 6408 4536
rect 4959 4499 5017 4505
rect 4522 4468 4528 4480
rect 3568 4440 4528 4468
rect 3568 4428 3574 4440
rect 4522 4428 4528 4440
rect 4580 4468 4586 4480
rect 5442 4468 5448 4480
rect 4580 4440 5448 4468
rect 4580 4428 4586 4440
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 5626 4468 5632 4480
rect 5583 4440 5632 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 1104 4378 6968 4400
rect 1104 4326 2376 4378
rect 2428 4326 2440 4378
rect 2492 4326 2504 4378
rect 2556 4326 2568 4378
rect 2620 4326 2632 4378
rect 2684 4326 3802 4378
rect 3854 4326 3866 4378
rect 3918 4326 3930 4378
rect 3982 4326 3994 4378
rect 4046 4326 4058 4378
rect 4110 4326 5228 4378
rect 5280 4326 5292 4378
rect 5344 4326 5356 4378
rect 5408 4326 5420 4378
rect 5472 4326 5484 4378
rect 5536 4326 6654 4378
rect 6706 4326 6718 4378
rect 6770 4326 6782 4378
rect 6834 4326 6846 4378
rect 6898 4326 6910 4378
rect 6962 4326 6968 4378
rect 1104 4304 6968 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 3660 4236 4292 4264
rect 3660 4224 3666 4236
rect 4264 4196 4292 4236
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4433 4267 4491 4273
rect 4433 4264 4445 4267
rect 4396 4236 4445 4264
rect 4396 4224 4402 4236
rect 4433 4233 4445 4236
rect 4479 4233 4491 4267
rect 4433 4227 4491 4233
rect 4724 4236 5120 4264
rect 4724 4196 4752 4236
rect 4982 4196 4988 4208
rect 4264 4168 4752 4196
rect 4816 4168 4988 4196
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 3712 4060 3740 4091
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4028 4100 4353 4128
rect 4028 4088 4034 4100
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4816 4128 4844 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 5092 4137 5120 4236
rect 5718 4224 5724 4276
rect 5776 4224 5782 4276
rect 5905 4267 5963 4273
rect 5905 4233 5917 4267
rect 5951 4264 5963 4267
rect 5994 4264 6000 4276
rect 5951 4236 6000 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 5736 4196 5764 4224
rect 5736 4168 6040 4196
rect 4663 4100 4844 4128
rect 4893 4131 4951 4137
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4893 4097 4905 4131
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5350 4128 5356 4140
rect 5307 4100 5356 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 4062 4060 4068 4072
rect 3712 4032 4068 4060
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4060 4307 4063
rect 4540 4060 4568 4088
rect 4295 4032 4568 4060
rect 4908 4060 4936 4091
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 6012 4137 6040 4168
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 5997 4131 6055 4137
rect 5767 4100 5856 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 5644 4060 5672 4088
rect 5828 4072 5856 4100
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6362 4128 6368 4140
rect 6227 4100 6368 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 4908 4032 5672 4060
rect 4295 4029 4307 4032
rect 4249 4023 4307 4029
rect 5810 4020 5816 4072
rect 5868 4020 5874 4072
rect 3881 3995 3939 4001
rect 3881 3961 3893 3995
rect 3927 3992 3939 3995
rect 4338 3992 4344 4004
rect 3927 3964 4344 3992
rect 3927 3961 3939 3964
rect 3881 3955 3939 3961
rect 4338 3952 4344 3964
rect 4396 3952 4402 4004
rect 5074 3952 5080 4004
rect 5132 3992 5138 4004
rect 5997 3995 6055 4001
rect 5997 3992 6009 3995
rect 5132 3964 6009 3992
rect 5132 3952 5138 3964
rect 5997 3961 6009 3964
rect 6043 3961 6055 3995
rect 5997 3955 6055 3961
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4246 3884 4252 3936
rect 4304 3884 4310 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 6546 3924 6552 3936
rect 5408 3896 6552 3924
rect 5408 3884 5414 3896
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 1104 3834 6808 3856
rect 1104 3782 1663 3834
rect 1715 3782 1727 3834
rect 1779 3782 1791 3834
rect 1843 3782 1855 3834
rect 1907 3782 1919 3834
rect 1971 3782 3089 3834
rect 3141 3782 3153 3834
rect 3205 3782 3217 3834
rect 3269 3782 3281 3834
rect 3333 3782 3345 3834
rect 3397 3782 4515 3834
rect 4567 3782 4579 3834
rect 4631 3782 4643 3834
rect 4695 3782 4707 3834
rect 4759 3782 4771 3834
rect 4823 3782 5941 3834
rect 5993 3782 6005 3834
rect 6057 3782 6069 3834
rect 6121 3782 6133 3834
rect 6185 3782 6197 3834
rect 6249 3782 6808 3834
rect 1104 3760 6808 3782
rect 3970 3680 3976 3732
rect 4028 3680 4034 3732
rect 4154 3680 4160 3732
rect 4212 3680 4218 3732
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 4488 3692 4629 3720
rect 4488 3680 4494 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 4617 3683 4675 3689
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5500 3692 5917 3720
rect 5500 3680 5506 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 5994 3680 6000 3732
rect 6052 3680 6058 3732
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6457 3723 6515 3729
rect 6457 3720 6469 3723
rect 6328 3692 6469 3720
rect 6328 3680 6334 3692
rect 6457 3689 6469 3692
rect 6503 3689 6515 3723
rect 6457 3683 6515 3689
rect 3988 3584 4016 3680
rect 2792 3556 4016 3584
rect 2792 3525 2820 3556
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1581 3451 1639 3457
rect 1581 3448 1593 3451
rect 992 3420 1593 3448
rect 992 3408 998 3420
rect 1581 3417 1593 3420
rect 1627 3417 1639 3451
rect 3804 3448 3832 3479
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 4172 3516 4200 3680
rect 4448 3624 6224 3652
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 4172 3488 4353 3516
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4448 3448 4476 3624
rect 6196 3596 6224 3624
rect 4522 3544 4528 3596
rect 4580 3544 4586 3596
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 4816 3556 6101 3584
rect 4540 3516 4568 3544
rect 4816 3525 4844 3556
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4540 3488 4813 3516
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5276 3525 5304 3556
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 6178 3544 6184 3596
rect 6236 3544 6242 3596
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5626 3516 5632 3528
rect 5491 3488 5632 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 5721 3479 5779 3485
rect 6104 3488 6285 3516
rect 3804 3420 4476 3448
rect 4908 3448 4936 3476
rect 5736 3448 5764 3479
rect 5997 3451 6055 3457
rect 5997 3448 6009 3451
rect 4908 3420 6009 3448
rect 1581 3411 1639 3417
rect 5997 3417 6009 3420
rect 6043 3417 6055 3451
rect 5997 3411 6055 3417
rect 6104 3392 6132 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4154 3380 4160 3392
rect 4019 3352 4160 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4249 3383 4307 3389
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 4338 3380 4344 3392
rect 4295 3352 4344 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4525 3383 4583 3389
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 5350 3380 5356 3392
rect 4571 3352 5356 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 6086 3340 6092 3392
rect 6144 3340 6150 3392
rect 1104 3290 6968 3312
rect 1104 3238 2376 3290
rect 2428 3238 2440 3290
rect 2492 3238 2504 3290
rect 2556 3238 2568 3290
rect 2620 3238 2632 3290
rect 2684 3238 3802 3290
rect 3854 3238 3866 3290
rect 3918 3238 3930 3290
rect 3982 3238 3994 3290
rect 4046 3238 4058 3290
rect 4110 3238 5228 3290
rect 5280 3238 5292 3290
rect 5344 3238 5356 3290
rect 5408 3238 5420 3290
rect 5472 3238 5484 3290
rect 5536 3238 6654 3290
rect 6706 3238 6718 3290
rect 6770 3238 6782 3290
rect 6834 3238 6846 3290
rect 6898 3238 6910 3290
rect 6962 3238 6968 3290
rect 1104 3216 6968 3238
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 4890 3176 4896 3188
rect 4847 3148 4896 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 4982 3136 4988 3188
rect 5040 3176 5046 3188
rect 5258 3176 5264 3188
rect 5040 3148 5264 3176
rect 5040 3136 5046 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 5626 3176 5632 3188
rect 5491 3148 5632 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 6380 3108 6408 3136
rect 5000 3080 6408 3108
rect 4246 3000 4252 3052
rect 4304 3000 4310 3052
rect 5000 3049 5028 3080
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 4338 2932 4344 2984
rect 4396 2932 4402 2984
rect 4356 2836 4384 2932
rect 4433 2907 4491 2913
rect 4433 2873 4445 2907
rect 4479 2904 4491 2907
rect 4540 2904 4568 3003
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 5092 2972 5120 3003
rect 5166 3000 5172 3052
rect 5224 3000 5230 3052
rect 5350 3000 5356 3052
rect 5408 3000 5414 3052
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5500 3012 5641 3040
rect 5500 3000 5506 3012
rect 5629 3009 5641 3012
rect 5675 3040 5687 3043
rect 5810 3040 5816 3052
rect 5675 3012 5816 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 5920 2972 5948 3003
rect 6086 3000 6092 3052
rect 6144 3000 6150 3052
rect 4663 2944 5120 2972
rect 5368 2944 5948 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 5074 2904 5080 2916
rect 4479 2876 5080 2904
rect 4479 2873 4491 2876
rect 4433 2867 4491 2873
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 5368 2913 5396 2944
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2873 5411 2907
rect 5353 2867 5411 2873
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6104 2904 6132 3000
rect 5868 2876 6132 2904
rect 5868 2864 5874 2876
rect 5442 2836 5448 2848
rect 4356 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 1104 2746 6808 2768
rect 1104 2694 1663 2746
rect 1715 2694 1727 2746
rect 1779 2694 1791 2746
rect 1843 2694 1855 2746
rect 1907 2694 1919 2746
rect 1971 2694 3089 2746
rect 3141 2694 3153 2746
rect 3205 2694 3217 2746
rect 3269 2694 3281 2746
rect 3333 2694 3345 2746
rect 3397 2694 4515 2746
rect 4567 2694 4579 2746
rect 4631 2694 4643 2746
rect 4695 2694 4707 2746
rect 4759 2694 4771 2746
rect 4823 2694 5941 2746
rect 5993 2694 6005 2746
rect 6057 2694 6069 2746
rect 6121 2694 6133 2746
rect 6185 2694 6197 2746
rect 6249 2694 6808 2746
rect 1104 2672 6808 2694
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5166 2632 5172 2644
rect 4939 2604 5172 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5258 2592 5264 2644
rect 5316 2632 5322 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5316 2604 6009 2632
rect 5316 2592 5322 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 4985 2567 5043 2573
rect 4985 2533 4997 2567
rect 5031 2564 5043 2567
rect 5350 2564 5356 2576
rect 5031 2536 5356 2564
rect 5031 2533 5043 2536
rect 4985 2527 5043 2533
rect 5350 2524 5356 2536
rect 5408 2564 5414 2576
rect 5629 2567 5687 2573
rect 5629 2564 5641 2567
rect 5408 2536 5641 2564
rect 5408 2524 5414 2536
rect 5629 2533 5641 2536
rect 5675 2533 5687 2567
rect 5629 2527 5687 2533
rect 5810 2524 5816 2576
rect 5868 2524 5874 2576
rect 4172 2468 4844 2496
rect 4172 2440 4200 2468
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2774 2428 2780 2440
rect 2731 2400 2780 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4632 2400 4721 2428
rect 1578 2320 1584 2372
rect 1636 2320 1642 2372
rect 4632 2292 4660 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4816 2360 4844 2468
rect 4890 2456 4896 2508
rect 4948 2496 4954 2508
rect 5828 2496 5856 2524
rect 4948 2468 5212 2496
rect 4948 2456 4954 2468
rect 5184 2437 5212 2468
rect 5276 2468 5856 2496
rect 5276 2437 5304 2468
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 5276 2360 5304 2391
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2428 5595 2431
rect 5626 2428 5632 2440
rect 5583 2400 5632 2428
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 4816 2332 5304 2360
rect 5353 2363 5411 2369
rect 5353 2329 5365 2363
rect 5399 2360 5411 2363
rect 5828 2360 5856 2391
rect 5399 2332 5856 2360
rect 5399 2329 5411 2332
rect 5353 2323 5411 2329
rect 6178 2320 6184 2372
rect 6236 2320 6242 2372
rect 6196 2292 6224 2320
rect 4632 2264 6224 2292
rect 1104 2202 6968 2224
rect 1104 2150 2376 2202
rect 2428 2150 2440 2202
rect 2492 2150 2504 2202
rect 2556 2150 2568 2202
rect 2620 2150 2632 2202
rect 2684 2150 3802 2202
rect 3854 2150 3866 2202
rect 3918 2150 3930 2202
rect 3982 2150 3994 2202
rect 4046 2150 4058 2202
rect 4110 2150 5228 2202
rect 5280 2150 5292 2202
rect 5344 2150 5356 2202
rect 5408 2150 5420 2202
rect 5472 2150 5484 2202
rect 5536 2150 6654 2202
rect 6706 2150 6718 2202
rect 6770 2150 6782 2202
rect 6834 2150 6846 2202
rect 6898 2150 6910 2202
rect 6962 2150 6968 2202
rect 1104 2128 6968 2150
rect 5074 2048 5080 2100
rect 5132 2088 5138 2100
rect 5626 2088 5632 2100
rect 5132 2060 5632 2088
rect 5132 2048 5138 2060
rect 5626 2048 5632 2060
rect 5684 2048 5690 2100
<< via1 >>
rect 4988 5720 5040 5772
rect 6276 5720 6328 5772
rect 3516 5584 3568 5636
rect 4804 5516 4856 5568
rect 5632 5516 5684 5568
rect 5724 5516 5776 5568
rect 2376 5414 2428 5466
rect 2440 5414 2492 5466
rect 2504 5414 2556 5466
rect 2568 5414 2620 5466
rect 2632 5414 2684 5466
rect 3802 5414 3854 5466
rect 3866 5414 3918 5466
rect 3930 5414 3982 5466
rect 3994 5414 4046 5466
rect 4058 5414 4110 5466
rect 5228 5414 5280 5466
rect 5292 5414 5344 5466
rect 5356 5414 5408 5466
rect 5420 5414 5472 5466
rect 5484 5414 5536 5466
rect 6654 5414 6706 5466
rect 6718 5414 6770 5466
rect 6782 5414 6834 5466
rect 6846 5414 6898 5466
rect 6910 5414 6962 5466
rect 3056 5312 3108 5364
rect 3240 5312 3292 5364
rect 3424 5312 3476 5364
rect 3516 5244 3568 5296
rect 940 5108 992 5160
rect 3332 5176 3384 5228
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 6368 5312 6420 5364
rect 4712 5244 4764 5296
rect 5540 5244 5592 5296
rect 4436 5176 4488 5228
rect 4896 5176 4948 5228
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 6460 5244 6512 5296
rect 5172 5176 5224 5185
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 4712 5040 4764 5092
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 6552 5176 6604 5228
rect 5356 5040 5408 5092
rect 3516 4972 3568 5024
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 4160 4972 4212 4981
rect 4252 4972 4304 5024
rect 5264 4972 5316 5024
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 1663 4870 1715 4922
rect 1727 4870 1779 4922
rect 1791 4870 1843 4922
rect 1855 4870 1907 4922
rect 1919 4870 1971 4922
rect 3089 4870 3141 4922
rect 3153 4870 3205 4922
rect 3217 4870 3269 4922
rect 3281 4870 3333 4922
rect 3345 4870 3397 4922
rect 4515 4870 4567 4922
rect 4579 4870 4631 4922
rect 4643 4870 4695 4922
rect 4707 4870 4759 4922
rect 4771 4870 4823 4922
rect 5941 4870 5993 4922
rect 6005 4870 6057 4922
rect 6069 4870 6121 4922
rect 6133 4870 6185 4922
rect 6197 4870 6249 4922
rect 3792 4768 3844 4820
rect 4896 4768 4948 4820
rect 5356 4768 5408 4820
rect 5448 4768 5500 4820
rect 2780 4700 2832 4752
rect 3332 4700 3384 4752
rect 4068 4700 4120 4752
rect 4344 4700 4396 4752
rect 2964 4564 3016 4616
rect 3332 4564 3384 4616
rect 3700 4564 3752 4616
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 2780 4496 2832 4548
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 3424 4428 3476 4480
rect 3516 4428 3568 4480
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 5264 4632 5316 4684
rect 4804 4564 4856 4573
rect 5632 4564 5684 4616
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6368 4564 6420 4616
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 4528 4428 4580 4480
rect 5448 4428 5500 4480
rect 5632 4428 5684 4480
rect 2376 4326 2428 4378
rect 2440 4326 2492 4378
rect 2504 4326 2556 4378
rect 2568 4326 2620 4378
rect 2632 4326 2684 4378
rect 3802 4326 3854 4378
rect 3866 4326 3918 4378
rect 3930 4326 3982 4378
rect 3994 4326 4046 4378
rect 4058 4326 4110 4378
rect 5228 4326 5280 4378
rect 5292 4326 5344 4378
rect 5356 4326 5408 4378
rect 5420 4326 5472 4378
rect 5484 4326 5536 4378
rect 6654 4326 6706 4378
rect 6718 4326 6770 4378
rect 6782 4326 6834 4378
rect 6846 4326 6898 4378
rect 6910 4326 6962 4378
rect 3608 4224 3660 4276
rect 4344 4224 4396 4276
rect 3976 4088 4028 4140
rect 4528 4088 4580 4140
rect 4988 4156 5040 4208
rect 5724 4224 5776 4276
rect 6000 4224 6052 4276
rect 4068 4020 4120 4072
rect 5356 4088 5408 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 5632 4088 5684 4140
rect 6368 4088 6420 4140
rect 5816 4020 5868 4072
rect 4344 3952 4396 4004
rect 5080 3952 5132 4004
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 4252 3927 4304 3936
rect 4252 3893 4261 3927
rect 4261 3893 4295 3927
rect 4295 3893 4304 3927
rect 4252 3884 4304 3893
rect 5356 3884 5408 3936
rect 6552 3884 6604 3936
rect 1663 3782 1715 3834
rect 1727 3782 1779 3834
rect 1791 3782 1843 3834
rect 1855 3782 1907 3834
rect 1919 3782 1971 3834
rect 3089 3782 3141 3834
rect 3153 3782 3205 3834
rect 3217 3782 3269 3834
rect 3281 3782 3333 3834
rect 3345 3782 3397 3834
rect 4515 3782 4567 3834
rect 4579 3782 4631 3834
rect 4643 3782 4695 3834
rect 4707 3782 4759 3834
rect 4771 3782 4823 3834
rect 5941 3782 5993 3834
rect 6005 3782 6057 3834
rect 6069 3782 6121 3834
rect 6133 3782 6185 3834
rect 6197 3782 6249 3834
rect 3976 3680 4028 3732
rect 4160 3680 4212 3732
rect 4436 3680 4488 3732
rect 5448 3680 5500 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 6276 3680 6328 3732
rect 940 3408 992 3460
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4528 3544 4580 3596
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 6184 3544 6236 3596
rect 5632 3476 5684 3528
rect 4160 3340 4212 3392
rect 4344 3340 4396 3392
rect 5356 3340 5408 3392
rect 6092 3340 6144 3392
rect 2376 3238 2428 3290
rect 2440 3238 2492 3290
rect 2504 3238 2556 3290
rect 2568 3238 2620 3290
rect 2632 3238 2684 3290
rect 3802 3238 3854 3290
rect 3866 3238 3918 3290
rect 3930 3238 3982 3290
rect 3994 3238 4046 3290
rect 4058 3238 4110 3290
rect 5228 3238 5280 3290
rect 5292 3238 5344 3290
rect 5356 3238 5408 3290
rect 5420 3238 5472 3290
rect 5484 3238 5536 3290
rect 6654 3238 6706 3290
rect 6718 3238 6770 3290
rect 6782 3238 6834 3290
rect 6846 3238 6898 3290
rect 6910 3238 6962 3290
rect 4896 3136 4948 3188
rect 4988 3136 5040 3188
rect 5264 3136 5316 3188
rect 5632 3136 5684 3188
rect 6368 3136 6420 3188
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 4344 2932 4396 2984
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 5448 3000 5500 3052
rect 5816 3000 5868 3052
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 5080 2864 5132 2916
rect 5816 2864 5868 2916
rect 5448 2796 5500 2848
rect 1663 2694 1715 2746
rect 1727 2694 1779 2746
rect 1791 2694 1843 2746
rect 1855 2694 1907 2746
rect 1919 2694 1971 2746
rect 3089 2694 3141 2746
rect 3153 2694 3205 2746
rect 3217 2694 3269 2746
rect 3281 2694 3333 2746
rect 3345 2694 3397 2746
rect 4515 2694 4567 2746
rect 4579 2694 4631 2746
rect 4643 2694 4695 2746
rect 4707 2694 4759 2746
rect 4771 2694 4823 2746
rect 5941 2694 5993 2746
rect 6005 2694 6057 2746
rect 6069 2694 6121 2746
rect 6133 2694 6185 2746
rect 6197 2694 6249 2746
rect 5172 2592 5224 2644
rect 5264 2592 5316 2644
rect 5356 2524 5408 2576
rect 5816 2524 5868 2576
rect 2780 2388 2832 2440
rect 4160 2388 4212 2440
rect 1584 2363 1636 2372
rect 1584 2329 1593 2363
rect 1593 2329 1627 2363
rect 1627 2329 1636 2363
rect 1584 2320 1636 2329
rect 4896 2456 4948 2508
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 5632 2388 5684 2440
rect 6184 2320 6236 2372
rect 2376 2150 2428 2202
rect 2440 2150 2492 2202
rect 2504 2150 2556 2202
rect 2568 2150 2620 2202
rect 2632 2150 2684 2202
rect 3802 2150 3854 2202
rect 3866 2150 3918 2202
rect 3930 2150 3982 2202
rect 3994 2150 4046 2202
rect 4058 2150 4110 2202
rect 5228 2150 5280 2202
rect 5292 2150 5344 2202
rect 5356 2150 5408 2202
rect 5420 2150 5472 2202
rect 5484 2150 5536 2202
rect 6654 2150 6706 2202
rect 6718 2150 6770 2202
rect 6782 2150 6834 2202
rect 6846 2150 6898 2202
rect 6910 2150 6962 2202
rect 5080 2048 5132 2100
rect 5632 2048 5684 2100
<< metal2 >>
rect 3790 6080 3846 6089
rect 3712 6038 3790 6066
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 3054 5808 3110 5817
rect 3054 5743 3110 5752
rect 2376 5468 2684 5477
rect 2376 5466 2382 5468
rect 2438 5466 2462 5468
rect 2518 5466 2542 5468
rect 2598 5466 2622 5468
rect 2678 5466 2684 5468
rect 2438 5414 2440 5466
rect 2620 5414 2622 5466
rect 2376 5412 2382 5414
rect 2438 5412 2462 5414
rect 2518 5412 2542 5414
rect 2598 5412 2622 5414
rect 2678 5412 2684 5414
rect 2376 5403 2684 5412
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 5001 980 5102
rect 938 4992 994 5001
rect 938 4927 994 4936
rect 1663 4924 1971 4933
rect 1663 4922 1669 4924
rect 1725 4922 1749 4924
rect 1805 4922 1829 4924
rect 1885 4922 1909 4924
rect 1965 4922 1971 4924
rect 1725 4870 1727 4922
rect 1907 4870 1909 4922
rect 1663 4868 1669 4870
rect 1725 4868 1749 4870
rect 1805 4868 1829 4870
rect 1885 4868 1909 4870
rect 1965 4868 1971 4870
rect 1663 4859 1971 4868
rect 2792 4758 2820 5743
rect 3068 5370 3096 5743
rect 3330 5672 3386 5681
rect 3252 5630 3330 5658
rect 3252 5370 3280 5630
rect 3330 5607 3386 5616
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3344 5137 3372 5170
rect 3330 5128 3386 5137
rect 3330 5063 3386 5072
rect 3089 4924 3397 4933
rect 3089 4922 3095 4924
rect 3151 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3397 4924
rect 3151 4870 3153 4922
rect 3333 4870 3335 4922
rect 3089 4868 3095 4870
rect 3151 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3397 4870
rect 3089 4859 3397 4868
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3344 4622 3372 4694
rect 2964 4616 3016 4622
rect 2962 4584 2964 4593
rect 3332 4616 3384 4622
rect 3016 4584 3018 4593
rect 2780 4548 2832 4554
rect 3332 4558 3384 4564
rect 2962 4519 3018 4528
rect 2780 4490 2832 4496
rect 2376 4380 2684 4389
rect 2376 4378 2382 4380
rect 2438 4378 2462 4380
rect 2518 4378 2542 4380
rect 2598 4378 2622 4380
rect 2678 4378 2684 4380
rect 2438 4326 2440 4378
rect 2620 4326 2622 4378
rect 2376 4324 2382 4326
rect 2438 4324 2462 4326
rect 2518 4324 2542 4326
rect 2598 4324 2622 4326
rect 2678 4324 2684 4326
rect 2376 4315 2684 4324
rect 1663 3836 1971 3845
rect 1663 3834 1669 3836
rect 1725 3834 1749 3836
rect 1805 3834 1829 3836
rect 1885 3834 1909 3836
rect 1965 3834 1971 3836
rect 1725 3782 1727 3834
rect 1907 3782 1909 3834
rect 1663 3780 1669 3782
rect 1725 3780 1749 3782
rect 1805 3780 1829 3782
rect 1885 3780 1909 3782
rect 1965 3780 1971 3782
rect 1663 3771 1971 3780
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3097 980 3402
rect 2376 3292 2684 3301
rect 2376 3290 2382 3292
rect 2438 3290 2462 3292
rect 2518 3290 2542 3292
rect 2598 3290 2622 3292
rect 2678 3290 2684 3292
rect 2438 3238 2440 3290
rect 2620 3238 2622 3290
rect 2376 3236 2382 3238
rect 2438 3236 2462 3238
rect 2518 3236 2542 3238
rect 2598 3236 2622 3238
rect 2678 3236 2684 3238
rect 2376 3227 2684 3236
rect 938 3088 994 3097
rect 938 3023 994 3032
rect 1663 2748 1971 2757
rect 1663 2746 1669 2748
rect 1725 2746 1749 2748
rect 1805 2746 1829 2748
rect 1885 2746 1909 2748
rect 1965 2746 1971 2748
rect 1725 2694 1727 2746
rect 1907 2694 1909 2746
rect 1663 2692 1669 2694
rect 1725 2692 1749 2694
rect 1805 2692 1829 2694
rect 1885 2692 1909 2694
rect 1965 2692 1971 2694
rect 1663 2683 1971 2692
rect 2792 2446 2820 4490
rect 3436 4486 3464 5306
rect 3528 5302 3556 5578
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3606 5264 3662 5273
rect 3606 5199 3662 5208
rect 3620 5030 3648 5199
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3528 4486 3556 4966
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3068 4049 3096 4422
rect 3620 4282 3648 4966
rect 3712 4622 3740 6038
rect 3790 6015 3846 6024
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 3802 5468 4110 5477
rect 3802 5466 3808 5468
rect 3864 5466 3888 5468
rect 3944 5466 3968 5468
rect 4024 5466 4048 5468
rect 4104 5466 4110 5468
rect 3864 5414 3866 5466
rect 4046 5414 4048 5466
rect 3802 5412 3808 5414
rect 3864 5412 3888 5414
rect 3944 5412 3968 5414
rect 4024 5412 4048 5414
rect 4104 5412 4110 5414
rect 3802 5403 4110 5412
rect 4356 5358 4752 5386
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3896 5114 3924 5170
rect 3896 5086 4292 5114
rect 4264 5030 4292 5086
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3804 4622 3832 4762
rect 4068 4752 4120 4758
rect 4066 4720 4068 4729
rect 4120 4720 4122 4729
rect 4066 4655 4122 4664
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3802 4380 4110 4389
rect 3802 4378 3808 4380
rect 3864 4378 3888 4380
rect 3944 4378 3968 4380
rect 4024 4378 4048 4380
rect 4104 4378 4110 4380
rect 3864 4326 3866 4378
rect 4046 4326 4048 4378
rect 3802 4324 3808 4326
rect 3864 4324 3888 4326
rect 3944 4324 3968 4326
rect 4024 4324 4048 4326
rect 4104 4324 4110 4326
rect 3802 4315 4110 4324
rect 3608 4276 3660 4282
rect 4172 4264 4200 4966
rect 4356 4758 4384 5358
rect 4724 5302 4752 5358
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4344 4752 4396 4758
rect 3608 4218 3660 4224
rect 3988 4236 4200 4264
rect 4264 4700 4344 4706
rect 4264 4694 4396 4700
rect 4264 4678 4384 4694
rect 3988 4146 4016 4236
rect 4066 4176 4122 4185
rect 3976 4140 4028 4146
rect 4122 4134 4200 4162
rect 4066 4111 4122 4120
rect 3976 4082 4028 4088
rect 4068 4072 4120 4078
rect 3054 4040 3110 4049
rect 4068 4014 4120 4020
rect 3054 3975 3110 3984
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3089 3836 3397 3845
rect 3089 3834 3095 3836
rect 3151 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3397 3836
rect 3151 3782 3153 3834
rect 3333 3782 3335 3834
rect 3089 3780 3095 3782
rect 3151 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3397 3782
rect 3089 3771 3397 3780
rect 3988 3738 4016 3878
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3641 4108 4014
rect 4172 3738 4200 4134
rect 4264 3942 4292 4678
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4356 4282 4384 4558
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4066 3632 4122 3641
rect 4356 3618 4384 3946
rect 4448 3738 4476 5170
rect 4816 5114 4844 5510
rect 5000 5234 5028 5714
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5228 5468 5536 5477
rect 5228 5466 5234 5468
rect 5290 5466 5314 5468
rect 5370 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5536 5468
rect 5290 5414 5292 5466
rect 5472 5414 5474 5466
rect 5228 5412 5234 5414
rect 5290 5412 5314 5414
rect 5370 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5536 5414
rect 5228 5403 5536 5412
rect 5540 5296 5592 5302
rect 5368 5273 5540 5284
rect 5354 5264 5540 5273
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5172 5228 5224 5234
rect 5410 5256 5540 5264
rect 5540 5238 5592 5244
rect 5354 5199 5410 5208
rect 5172 5170 5224 5176
rect 4724 5098 4844 5114
rect 4712 5092 4844 5098
rect 4764 5086 4844 5092
rect 4712 5034 4764 5040
rect 4515 4924 4823 4933
rect 4515 4922 4521 4924
rect 4577 4922 4601 4924
rect 4657 4922 4681 4924
rect 4737 4922 4761 4924
rect 4817 4922 4823 4924
rect 4577 4870 4579 4922
rect 4759 4870 4761 4922
rect 4515 4868 4521 4870
rect 4577 4868 4601 4870
rect 4657 4868 4681 4870
rect 4737 4868 4761 4870
rect 4817 4868 4823 4870
rect 4515 4859 4823 4868
rect 4908 4826 4936 5170
rect 5080 5160 5132 5166
rect 4986 5128 5042 5137
rect 5080 5102 5132 5108
rect 4986 5063 5042 5072
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4616 4856 4622
rect 4856 4576 4936 4604
rect 4804 4558 4856 4564
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4540 4146 4568 4422
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4908 3890 4936 4576
rect 5000 4214 5028 5063
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5092 4010 5120 5102
rect 5184 4672 5212 5170
rect 5540 5160 5592 5166
rect 5446 5128 5502 5137
rect 5356 5092 5408 5098
rect 5540 5102 5592 5108
rect 5446 5063 5502 5072
rect 5356 5034 5408 5040
rect 5264 5024 5316 5030
rect 5262 4992 5264 5001
rect 5316 4992 5318 5001
rect 5262 4927 5318 4936
rect 5368 4826 5396 5034
rect 5460 5030 5488 5063
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4826 5488 4966
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5264 4684 5316 4690
rect 5184 4644 5264 4672
rect 5264 4626 5316 4632
rect 5448 4480 5500 4486
rect 5552 4468 5580 5102
rect 5644 4622 5672 5510
rect 5736 5273 5764 5510
rect 5722 5264 5778 5273
rect 5722 5199 5778 5208
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 6012 5012 6040 5170
rect 5736 4984 6040 5012
rect 5736 4740 5764 4984
rect 5941 4924 6249 4933
rect 5941 4922 5947 4924
rect 6003 4922 6027 4924
rect 6083 4922 6107 4924
rect 6163 4922 6187 4924
rect 6243 4922 6249 4924
rect 6003 4870 6005 4922
rect 6185 4870 6187 4922
rect 5941 4868 5947 4870
rect 6003 4868 6027 4870
rect 6083 4868 6107 4870
rect 6163 4868 6187 4870
rect 6243 4868 6249 4870
rect 5941 4859 6249 4868
rect 5736 4712 5856 4740
rect 5632 4616 5684 4622
rect 5684 4576 5764 4604
rect 5632 4558 5684 4564
rect 5500 4440 5580 4468
rect 5632 4480 5684 4486
rect 5448 4422 5500 4428
rect 5632 4422 5684 4428
rect 5228 4380 5536 4389
rect 5228 4378 5234 4380
rect 5290 4378 5314 4380
rect 5370 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5536 4380
rect 5290 4326 5292 4378
rect 5472 4326 5474 4378
rect 5228 4324 5234 4326
rect 5290 4324 5314 4326
rect 5370 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5536 4326
rect 5228 4315 5536 4324
rect 5644 4146 5672 4422
rect 5736 4282 5764 4576
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5368 3942 5396 4082
rect 5356 3936 5408 3942
rect 4908 3862 5120 3890
rect 5356 3878 5408 3884
rect 4515 3836 4823 3845
rect 4515 3834 4521 3836
rect 4577 3834 4601 3836
rect 4657 3834 4681 3836
rect 4737 3834 4761 3836
rect 4817 3834 4823 3836
rect 4577 3782 4579 3834
rect 4759 3782 4761 3834
rect 4515 3780 4521 3782
rect 4577 3780 4601 3782
rect 4657 3780 4681 3782
rect 4737 3780 4761 3782
rect 4817 3780 4823 3782
rect 4515 3771 4823 3780
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4356 3602 4568 3618
rect 4356 3596 4580 3602
rect 4356 3590 4528 3596
rect 4066 3567 4122 3576
rect 4528 3538 4580 3544
rect 5092 3534 5120 3862
rect 4068 3528 4120 3534
rect 4066 3496 4068 3505
rect 4896 3528 4948 3534
rect 4120 3496 4122 3505
rect 4896 3470 4948 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4066 3431 4122 3440
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 3802 3292 4110 3301
rect 3802 3290 3808 3292
rect 3864 3290 3888 3292
rect 3944 3290 3968 3292
rect 4024 3290 4048 3292
rect 4104 3290 4110 3292
rect 3864 3238 3866 3290
rect 4046 3238 4048 3290
rect 3802 3236 3808 3238
rect 3864 3236 3888 3238
rect 3944 3236 3968 3238
rect 4024 3236 4048 3238
rect 4104 3236 4110 3238
rect 3802 3227 4110 3236
rect 3089 2748 3397 2757
rect 3089 2746 3095 2748
rect 3151 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3397 2748
rect 3151 2694 3153 2746
rect 3333 2694 3335 2746
rect 3089 2692 3095 2694
rect 3151 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3397 2694
rect 3089 2683 3397 2692
rect 4172 2446 4200 3334
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4264 2774 4292 2994
rect 4356 2990 4384 3334
rect 4908 3194 4936 3470
rect 5000 3194 5028 3470
rect 5368 3398 5396 3878
rect 5460 3738 5488 4082
rect 5828 4078 5856 4712
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4282 6040 4558
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5816 4072 5868 4078
rect 5814 4040 5816 4049
rect 5868 4040 5870 4049
rect 5814 3975 5870 3984
rect 5941 3836 6249 3845
rect 5941 3834 5947 3836
rect 6003 3834 6027 3836
rect 6083 3834 6107 3836
rect 6163 3834 6187 3836
rect 6243 3834 6249 3836
rect 6003 3782 6005 3834
rect 6185 3782 6187 3834
rect 5941 3780 5947 3782
rect 6003 3780 6027 3782
rect 6083 3780 6107 3782
rect 6163 3780 6187 3782
rect 6243 3780 6249 3782
rect 5941 3771 6249 3780
rect 6288 3738 6316 5714
rect 6654 5468 6962 5477
rect 6654 5466 6660 5468
rect 6716 5466 6740 5468
rect 6796 5466 6820 5468
rect 6876 5466 6900 5468
rect 6956 5466 6962 5468
rect 6716 5414 6718 5466
rect 6898 5414 6900 5466
rect 6654 5412 6660 5414
rect 6716 5412 6740 5414
rect 6796 5412 6820 5414
rect 6876 5412 6900 5414
rect 6956 5412 6962 5414
rect 6654 5403 6962 5412
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6380 4622 6408 5306
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6472 4622 6500 5238
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6380 4146 6408 4558
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6564 3942 6592 5170
rect 6654 4380 6962 4389
rect 6654 4378 6660 4380
rect 6716 4378 6740 4380
rect 6796 4378 6820 4380
rect 6876 4378 6900 4380
rect 6956 4378 6962 4380
rect 6716 4326 6718 4378
rect 6898 4326 6900 4378
rect 6654 4324 6660 4326
rect 6716 4324 6740 4326
rect 6796 4324 6820 4326
rect 6876 4324 6900 4326
rect 6956 4324 6962 4326
rect 6654 4315 6962 4324
rect 6552 3936 6604 3942
rect 6366 3904 6422 3913
rect 6552 3878 6604 3884
rect 6366 3839 6422 3848
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6012 3618 6040 3674
rect 5920 3590 6040 3618
rect 6184 3596 6236 3602
rect 5632 3528 5684 3534
rect 5920 3482 5948 3590
rect 6184 3538 6236 3544
rect 5632 3470 5684 3476
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5228 3292 5536 3301
rect 5228 3290 5234 3292
rect 5290 3290 5314 3292
rect 5370 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5536 3292
rect 5290 3238 5292 3290
rect 5472 3238 5474 3290
rect 5228 3236 5234 3238
rect 5290 3236 5314 3238
rect 5370 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5536 3238
rect 5228 3227 5536 3236
rect 5644 3194 5672 3470
rect 5828 3454 5948 3482
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4894 2952 4950 2961
rect 4894 2887 4950 2896
rect 5080 2916 5132 2922
rect 4264 2746 4476 2774
rect 4448 2553 4476 2746
rect 4515 2748 4823 2757
rect 4515 2746 4521 2748
rect 4577 2746 4601 2748
rect 4657 2746 4681 2748
rect 4737 2746 4761 2748
rect 4817 2746 4823 2748
rect 4577 2694 4579 2746
rect 4759 2694 4761 2746
rect 4515 2692 4521 2694
rect 4577 2692 4601 2694
rect 4657 2692 4681 2694
rect 4737 2692 4761 2694
rect 4817 2692 4823 2694
rect 4515 2683 4823 2692
rect 4434 2544 4490 2553
rect 4908 2514 4936 2887
rect 5080 2858 5132 2864
rect 4434 2479 4490 2488
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1596 2045 1624 2314
rect 2376 2204 2684 2213
rect 2376 2202 2382 2204
rect 2438 2202 2462 2204
rect 2518 2202 2542 2204
rect 2598 2202 2622 2204
rect 2678 2202 2684 2204
rect 2438 2150 2440 2202
rect 2620 2150 2622 2202
rect 2376 2148 2382 2150
rect 2438 2148 2462 2150
rect 2518 2148 2542 2150
rect 2598 2148 2622 2150
rect 2678 2148 2684 2150
rect 2376 2139 2684 2148
rect 3802 2204 4110 2213
rect 3802 2202 3808 2204
rect 3864 2202 3888 2204
rect 3944 2202 3968 2204
rect 4024 2202 4048 2204
rect 4104 2202 4110 2204
rect 3864 2150 3866 2202
rect 4046 2150 4048 2202
rect 3802 2148 3808 2150
rect 3864 2148 3888 2150
rect 3944 2148 3968 2150
rect 4024 2148 4048 2150
rect 4104 2148 4110 2150
rect 3802 2139 4110 2148
rect 5092 2106 5120 2858
rect 5184 2650 5212 2994
rect 5276 2650 5304 3130
rect 5828 3058 5856 3454
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6104 3058 6132 3334
rect 6196 3097 6224 3538
rect 6380 3194 6408 3839
rect 6654 3292 6962 3301
rect 6654 3290 6660 3292
rect 6716 3290 6740 3292
rect 6796 3290 6820 3292
rect 6876 3290 6900 3292
rect 6956 3290 6962 3292
rect 6716 3238 6718 3290
rect 6898 3238 6900 3290
rect 6654 3236 6660 3238
rect 6716 3236 6740 3238
rect 6796 3236 6820 3238
rect 6876 3236 6900 3238
rect 6956 3236 6962 3238
rect 6654 3227 6962 3236
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6182 3088 6238 3097
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6092 3052 6144 3058
rect 6182 3023 6238 3032
rect 6092 2994 6144 3000
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5368 2582 5396 2994
rect 5460 2854 5488 2994
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 5460 2446 5488 2790
rect 5828 2582 5856 2858
rect 5941 2748 6249 2757
rect 5941 2746 5947 2748
rect 6003 2746 6027 2748
rect 6083 2746 6107 2748
rect 6163 2746 6187 2748
rect 6243 2746 6249 2748
rect 6003 2694 6005 2746
rect 6185 2694 6187 2746
rect 5941 2692 5947 2694
rect 6003 2692 6027 2694
rect 6083 2692 6107 2694
rect 6163 2692 6187 2694
rect 6243 2692 6249 2694
rect 5941 2683 6249 2692
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 6182 2408 6238 2417
rect 5228 2204 5536 2213
rect 5228 2202 5234 2204
rect 5290 2202 5314 2204
rect 5370 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5536 2204
rect 5290 2150 5292 2202
rect 5472 2150 5474 2202
rect 5228 2148 5234 2150
rect 5290 2148 5314 2150
rect 5370 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5536 2150
rect 5228 2139 5536 2148
rect 5644 2106 5672 2382
rect 6182 2343 6184 2352
rect 6236 2343 6238 2352
rect 6184 2314 6236 2320
rect 6654 2204 6962 2213
rect 6654 2202 6660 2204
rect 6716 2202 6740 2204
rect 6796 2202 6820 2204
rect 6876 2202 6900 2204
rect 6956 2202 6962 2204
rect 6716 2150 6718 2202
rect 6898 2150 6900 2202
rect 6654 2148 6660 2150
rect 6716 2148 6740 2150
rect 6796 2148 6820 2150
rect 6876 2148 6900 2150
rect 6956 2148 6962 2150
rect 6654 2139 6962 2148
rect 5080 2100 5132 2106
rect 1582 2036 1638 2045
rect 5080 2042 5132 2048
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 1582 1971 1638 1980
<< via2 >>
rect 2778 5752 2834 5808
rect 3054 5752 3110 5808
rect 2382 5466 2438 5468
rect 2462 5466 2518 5468
rect 2542 5466 2598 5468
rect 2622 5466 2678 5468
rect 2382 5414 2428 5466
rect 2428 5414 2438 5466
rect 2462 5414 2492 5466
rect 2492 5414 2504 5466
rect 2504 5414 2518 5466
rect 2542 5414 2556 5466
rect 2556 5414 2568 5466
rect 2568 5414 2598 5466
rect 2622 5414 2632 5466
rect 2632 5414 2678 5466
rect 2382 5412 2438 5414
rect 2462 5412 2518 5414
rect 2542 5412 2598 5414
rect 2622 5412 2678 5414
rect 938 4936 994 4992
rect 1669 4922 1725 4924
rect 1749 4922 1805 4924
rect 1829 4922 1885 4924
rect 1909 4922 1965 4924
rect 1669 4870 1715 4922
rect 1715 4870 1725 4922
rect 1749 4870 1779 4922
rect 1779 4870 1791 4922
rect 1791 4870 1805 4922
rect 1829 4870 1843 4922
rect 1843 4870 1855 4922
rect 1855 4870 1885 4922
rect 1909 4870 1919 4922
rect 1919 4870 1965 4922
rect 1669 4868 1725 4870
rect 1749 4868 1805 4870
rect 1829 4868 1885 4870
rect 1909 4868 1965 4870
rect 3330 5616 3386 5672
rect 3330 5072 3386 5128
rect 3095 4922 3151 4924
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3095 4870 3141 4922
rect 3141 4870 3151 4922
rect 3175 4870 3205 4922
rect 3205 4870 3217 4922
rect 3217 4870 3231 4922
rect 3255 4870 3269 4922
rect 3269 4870 3281 4922
rect 3281 4870 3311 4922
rect 3335 4870 3345 4922
rect 3345 4870 3391 4922
rect 3095 4868 3151 4870
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 2962 4564 2964 4584
rect 2964 4564 3016 4584
rect 3016 4564 3018 4584
rect 2962 4528 3018 4564
rect 2382 4378 2438 4380
rect 2462 4378 2518 4380
rect 2542 4378 2598 4380
rect 2622 4378 2678 4380
rect 2382 4326 2428 4378
rect 2428 4326 2438 4378
rect 2462 4326 2492 4378
rect 2492 4326 2504 4378
rect 2504 4326 2518 4378
rect 2542 4326 2556 4378
rect 2556 4326 2568 4378
rect 2568 4326 2598 4378
rect 2622 4326 2632 4378
rect 2632 4326 2678 4378
rect 2382 4324 2438 4326
rect 2462 4324 2518 4326
rect 2542 4324 2598 4326
rect 2622 4324 2678 4326
rect 1669 3834 1725 3836
rect 1749 3834 1805 3836
rect 1829 3834 1885 3836
rect 1909 3834 1965 3836
rect 1669 3782 1715 3834
rect 1715 3782 1725 3834
rect 1749 3782 1779 3834
rect 1779 3782 1791 3834
rect 1791 3782 1805 3834
rect 1829 3782 1843 3834
rect 1843 3782 1855 3834
rect 1855 3782 1885 3834
rect 1909 3782 1919 3834
rect 1919 3782 1965 3834
rect 1669 3780 1725 3782
rect 1749 3780 1805 3782
rect 1829 3780 1885 3782
rect 1909 3780 1965 3782
rect 2382 3290 2438 3292
rect 2462 3290 2518 3292
rect 2542 3290 2598 3292
rect 2622 3290 2678 3292
rect 2382 3238 2428 3290
rect 2428 3238 2438 3290
rect 2462 3238 2492 3290
rect 2492 3238 2504 3290
rect 2504 3238 2518 3290
rect 2542 3238 2556 3290
rect 2556 3238 2568 3290
rect 2568 3238 2598 3290
rect 2622 3238 2632 3290
rect 2632 3238 2678 3290
rect 2382 3236 2438 3238
rect 2462 3236 2518 3238
rect 2542 3236 2598 3238
rect 2622 3236 2678 3238
rect 938 3032 994 3088
rect 1669 2746 1725 2748
rect 1749 2746 1805 2748
rect 1829 2746 1885 2748
rect 1909 2746 1965 2748
rect 1669 2694 1715 2746
rect 1715 2694 1725 2746
rect 1749 2694 1779 2746
rect 1779 2694 1791 2746
rect 1791 2694 1805 2746
rect 1829 2694 1843 2746
rect 1843 2694 1855 2746
rect 1855 2694 1885 2746
rect 1909 2694 1919 2746
rect 1919 2694 1965 2746
rect 1669 2692 1725 2694
rect 1749 2692 1805 2694
rect 1829 2692 1885 2694
rect 1909 2692 1965 2694
rect 3606 5208 3662 5264
rect 3790 6024 3846 6080
rect 3808 5466 3864 5468
rect 3888 5466 3944 5468
rect 3968 5466 4024 5468
rect 4048 5466 4104 5468
rect 3808 5414 3854 5466
rect 3854 5414 3864 5466
rect 3888 5414 3918 5466
rect 3918 5414 3930 5466
rect 3930 5414 3944 5466
rect 3968 5414 3982 5466
rect 3982 5414 3994 5466
rect 3994 5414 4024 5466
rect 4048 5414 4058 5466
rect 4058 5414 4104 5466
rect 3808 5412 3864 5414
rect 3888 5412 3944 5414
rect 3968 5412 4024 5414
rect 4048 5412 4104 5414
rect 4066 4700 4068 4720
rect 4068 4700 4120 4720
rect 4120 4700 4122 4720
rect 4066 4664 4122 4700
rect 3808 4378 3864 4380
rect 3888 4378 3944 4380
rect 3968 4378 4024 4380
rect 4048 4378 4104 4380
rect 3808 4326 3854 4378
rect 3854 4326 3864 4378
rect 3888 4326 3918 4378
rect 3918 4326 3930 4378
rect 3930 4326 3944 4378
rect 3968 4326 3982 4378
rect 3982 4326 3994 4378
rect 3994 4326 4024 4378
rect 4048 4326 4058 4378
rect 4058 4326 4104 4378
rect 3808 4324 3864 4326
rect 3888 4324 3944 4326
rect 3968 4324 4024 4326
rect 4048 4324 4104 4326
rect 4066 4120 4122 4176
rect 3054 3984 3110 4040
rect 3095 3834 3151 3836
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3095 3782 3141 3834
rect 3141 3782 3151 3834
rect 3175 3782 3205 3834
rect 3205 3782 3217 3834
rect 3217 3782 3231 3834
rect 3255 3782 3269 3834
rect 3269 3782 3281 3834
rect 3281 3782 3311 3834
rect 3335 3782 3345 3834
rect 3345 3782 3391 3834
rect 3095 3780 3151 3782
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 4066 3576 4122 3632
rect 5234 5466 5290 5468
rect 5314 5466 5370 5468
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5234 5414 5280 5466
rect 5280 5414 5290 5466
rect 5314 5414 5344 5466
rect 5344 5414 5356 5466
rect 5356 5414 5370 5466
rect 5394 5414 5408 5466
rect 5408 5414 5420 5466
rect 5420 5414 5450 5466
rect 5474 5414 5484 5466
rect 5484 5414 5530 5466
rect 5234 5412 5290 5414
rect 5314 5412 5370 5414
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5354 5208 5410 5264
rect 4521 4922 4577 4924
rect 4601 4922 4657 4924
rect 4681 4922 4737 4924
rect 4761 4922 4817 4924
rect 4521 4870 4567 4922
rect 4567 4870 4577 4922
rect 4601 4870 4631 4922
rect 4631 4870 4643 4922
rect 4643 4870 4657 4922
rect 4681 4870 4695 4922
rect 4695 4870 4707 4922
rect 4707 4870 4737 4922
rect 4761 4870 4771 4922
rect 4771 4870 4817 4922
rect 4521 4868 4577 4870
rect 4601 4868 4657 4870
rect 4681 4868 4737 4870
rect 4761 4868 4817 4870
rect 4986 5072 5042 5128
rect 5446 5072 5502 5128
rect 5262 4972 5264 4992
rect 5264 4972 5316 4992
rect 5316 4972 5318 4992
rect 5262 4936 5318 4972
rect 5722 5208 5778 5264
rect 5947 4922 6003 4924
rect 6027 4922 6083 4924
rect 6107 4922 6163 4924
rect 6187 4922 6243 4924
rect 5947 4870 5993 4922
rect 5993 4870 6003 4922
rect 6027 4870 6057 4922
rect 6057 4870 6069 4922
rect 6069 4870 6083 4922
rect 6107 4870 6121 4922
rect 6121 4870 6133 4922
rect 6133 4870 6163 4922
rect 6187 4870 6197 4922
rect 6197 4870 6243 4922
rect 5947 4868 6003 4870
rect 6027 4868 6083 4870
rect 6107 4868 6163 4870
rect 6187 4868 6243 4870
rect 5234 4378 5290 4380
rect 5314 4378 5370 4380
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5234 4326 5280 4378
rect 5280 4326 5290 4378
rect 5314 4326 5344 4378
rect 5344 4326 5356 4378
rect 5356 4326 5370 4378
rect 5394 4326 5408 4378
rect 5408 4326 5420 4378
rect 5420 4326 5450 4378
rect 5474 4326 5484 4378
rect 5484 4326 5530 4378
rect 5234 4324 5290 4326
rect 5314 4324 5370 4326
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 4521 3834 4577 3836
rect 4601 3834 4657 3836
rect 4681 3834 4737 3836
rect 4761 3834 4817 3836
rect 4521 3782 4567 3834
rect 4567 3782 4577 3834
rect 4601 3782 4631 3834
rect 4631 3782 4643 3834
rect 4643 3782 4657 3834
rect 4681 3782 4695 3834
rect 4695 3782 4707 3834
rect 4707 3782 4737 3834
rect 4761 3782 4771 3834
rect 4771 3782 4817 3834
rect 4521 3780 4577 3782
rect 4601 3780 4657 3782
rect 4681 3780 4737 3782
rect 4761 3780 4817 3782
rect 4066 3476 4068 3496
rect 4068 3476 4120 3496
rect 4120 3476 4122 3496
rect 4066 3440 4122 3476
rect 3808 3290 3864 3292
rect 3888 3290 3944 3292
rect 3968 3290 4024 3292
rect 4048 3290 4104 3292
rect 3808 3238 3854 3290
rect 3854 3238 3864 3290
rect 3888 3238 3918 3290
rect 3918 3238 3930 3290
rect 3930 3238 3944 3290
rect 3968 3238 3982 3290
rect 3982 3238 3994 3290
rect 3994 3238 4024 3290
rect 4048 3238 4058 3290
rect 4058 3238 4104 3290
rect 3808 3236 3864 3238
rect 3888 3236 3944 3238
rect 3968 3236 4024 3238
rect 4048 3236 4104 3238
rect 3095 2746 3151 2748
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3095 2694 3141 2746
rect 3141 2694 3151 2746
rect 3175 2694 3205 2746
rect 3205 2694 3217 2746
rect 3217 2694 3231 2746
rect 3255 2694 3269 2746
rect 3269 2694 3281 2746
rect 3281 2694 3311 2746
rect 3335 2694 3345 2746
rect 3345 2694 3391 2746
rect 3095 2692 3151 2694
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 5814 4020 5816 4040
rect 5816 4020 5868 4040
rect 5868 4020 5870 4040
rect 5814 3984 5870 4020
rect 5947 3834 6003 3836
rect 6027 3834 6083 3836
rect 6107 3834 6163 3836
rect 6187 3834 6243 3836
rect 5947 3782 5993 3834
rect 5993 3782 6003 3834
rect 6027 3782 6057 3834
rect 6057 3782 6069 3834
rect 6069 3782 6083 3834
rect 6107 3782 6121 3834
rect 6121 3782 6133 3834
rect 6133 3782 6163 3834
rect 6187 3782 6197 3834
rect 6197 3782 6243 3834
rect 5947 3780 6003 3782
rect 6027 3780 6083 3782
rect 6107 3780 6163 3782
rect 6187 3780 6243 3782
rect 6660 5466 6716 5468
rect 6740 5466 6796 5468
rect 6820 5466 6876 5468
rect 6900 5466 6956 5468
rect 6660 5414 6706 5466
rect 6706 5414 6716 5466
rect 6740 5414 6770 5466
rect 6770 5414 6782 5466
rect 6782 5414 6796 5466
rect 6820 5414 6834 5466
rect 6834 5414 6846 5466
rect 6846 5414 6876 5466
rect 6900 5414 6910 5466
rect 6910 5414 6956 5466
rect 6660 5412 6716 5414
rect 6740 5412 6796 5414
rect 6820 5412 6876 5414
rect 6900 5412 6956 5414
rect 6660 4378 6716 4380
rect 6740 4378 6796 4380
rect 6820 4378 6876 4380
rect 6900 4378 6956 4380
rect 6660 4326 6706 4378
rect 6706 4326 6716 4378
rect 6740 4326 6770 4378
rect 6770 4326 6782 4378
rect 6782 4326 6796 4378
rect 6820 4326 6834 4378
rect 6834 4326 6846 4378
rect 6846 4326 6876 4378
rect 6900 4326 6910 4378
rect 6910 4326 6956 4378
rect 6660 4324 6716 4326
rect 6740 4324 6796 4326
rect 6820 4324 6876 4326
rect 6900 4324 6956 4326
rect 6366 3848 6422 3904
rect 5234 3290 5290 3292
rect 5314 3290 5370 3292
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5234 3238 5280 3290
rect 5280 3238 5290 3290
rect 5314 3238 5344 3290
rect 5344 3238 5356 3290
rect 5356 3238 5370 3290
rect 5394 3238 5408 3290
rect 5408 3238 5420 3290
rect 5420 3238 5450 3290
rect 5474 3238 5484 3290
rect 5484 3238 5530 3290
rect 5234 3236 5290 3238
rect 5314 3236 5370 3238
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 4894 2896 4950 2952
rect 4521 2746 4577 2748
rect 4601 2746 4657 2748
rect 4681 2746 4737 2748
rect 4761 2746 4817 2748
rect 4521 2694 4567 2746
rect 4567 2694 4577 2746
rect 4601 2694 4631 2746
rect 4631 2694 4643 2746
rect 4643 2694 4657 2746
rect 4681 2694 4695 2746
rect 4695 2694 4707 2746
rect 4707 2694 4737 2746
rect 4761 2694 4771 2746
rect 4771 2694 4817 2746
rect 4521 2692 4577 2694
rect 4601 2692 4657 2694
rect 4681 2692 4737 2694
rect 4761 2692 4817 2694
rect 4434 2488 4490 2544
rect 2382 2202 2438 2204
rect 2462 2202 2518 2204
rect 2542 2202 2598 2204
rect 2622 2202 2678 2204
rect 2382 2150 2428 2202
rect 2428 2150 2438 2202
rect 2462 2150 2492 2202
rect 2492 2150 2504 2202
rect 2504 2150 2518 2202
rect 2542 2150 2556 2202
rect 2556 2150 2568 2202
rect 2568 2150 2598 2202
rect 2622 2150 2632 2202
rect 2632 2150 2678 2202
rect 2382 2148 2438 2150
rect 2462 2148 2518 2150
rect 2542 2148 2598 2150
rect 2622 2148 2678 2150
rect 3808 2202 3864 2204
rect 3888 2202 3944 2204
rect 3968 2202 4024 2204
rect 4048 2202 4104 2204
rect 3808 2150 3854 2202
rect 3854 2150 3864 2202
rect 3888 2150 3918 2202
rect 3918 2150 3930 2202
rect 3930 2150 3944 2202
rect 3968 2150 3982 2202
rect 3982 2150 3994 2202
rect 3994 2150 4024 2202
rect 4048 2150 4058 2202
rect 4058 2150 4104 2202
rect 3808 2148 3864 2150
rect 3888 2148 3944 2150
rect 3968 2148 4024 2150
rect 4048 2148 4104 2150
rect 6660 3290 6716 3292
rect 6740 3290 6796 3292
rect 6820 3290 6876 3292
rect 6900 3290 6956 3292
rect 6660 3238 6706 3290
rect 6706 3238 6716 3290
rect 6740 3238 6770 3290
rect 6770 3238 6782 3290
rect 6782 3238 6796 3290
rect 6820 3238 6834 3290
rect 6834 3238 6846 3290
rect 6846 3238 6876 3290
rect 6900 3238 6910 3290
rect 6910 3238 6956 3290
rect 6660 3236 6716 3238
rect 6740 3236 6796 3238
rect 6820 3236 6876 3238
rect 6900 3236 6956 3238
rect 6182 3032 6238 3088
rect 5947 2746 6003 2748
rect 6027 2746 6083 2748
rect 6107 2746 6163 2748
rect 6187 2746 6243 2748
rect 5947 2694 5993 2746
rect 5993 2694 6003 2746
rect 6027 2694 6057 2746
rect 6057 2694 6069 2746
rect 6069 2694 6083 2746
rect 6107 2694 6121 2746
rect 6121 2694 6133 2746
rect 6133 2694 6163 2746
rect 6187 2694 6197 2746
rect 6197 2694 6243 2746
rect 5947 2692 6003 2694
rect 6027 2692 6083 2694
rect 6107 2692 6163 2694
rect 6187 2692 6243 2694
rect 5234 2202 5290 2204
rect 5314 2202 5370 2204
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5234 2150 5280 2202
rect 5280 2150 5290 2202
rect 5314 2150 5344 2202
rect 5344 2150 5356 2202
rect 5356 2150 5370 2202
rect 5394 2150 5408 2202
rect 5408 2150 5420 2202
rect 5420 2150 5450 2202
rect 5474 2150 5484 2202
rect 5484 2150 5530 2202
rect 5234 2148 5290 2150
rect 5314 2148 5370 2150
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 6182 2372 6238 2408
rect 6182 2352 6184 2372
rect 6184 2352 6236 2372
rect 6236 2352 6238 2372
rect 6660 2202 6716 2204
rect 6740 2202 6796 2204
rect 6820 2202 6876 2204
rect 6900 2202 6956 2204
rect 6660 2150 6706 2202
rect 6706 2150 6716 2202
rect 6740 2150 6770 2202
rect 6770 2150 6782 2202
rect 6782 2150 6796 2202
rect 6820 2150 6834 2202
rect 6834 2150 6846 2202
rect 6846 2150 6876 2202
rect 6900 2150 6910 2202
rect 6910 2150 6956 2202
rect 6660 2148 6716 2150
rect 6740 2148 6796 2150
rect 6820 2148 6876 2150
rect 6900 2148 6956 2150
rect 1582 1980 1638 2036
<< metal3 >>
rect 3785 6082 3851 6085
rect 7200 6082 8000 6112
rect 3785 6080 8000 6082
rect 3785 6024 3790 6080
rect 3846 6024 8000 6080
rect 3785 6022 8000 6024
rect 3785 6019 3851 6022
rect 7200 5992 8000 6022
rect 0 5810 800 5840
rect 2773 5810 2839 5813
rect 0 5808 2839 5810
rect 0 5752 2778 5808
rect 2834 5752 2839 5808
rect 0 5750 2839 5752
rect 0 5720 800 5750
rect 2773 5747 2839 5750
rect 3049 5810 3115 5813
rect 7200 5810 8000 5840
rect 3049 5808 8000 5810
rect 3049 5752 3054 5808
rect 3110 5752 8000 5808
rect 3049 5750 8000 5752
rect 3049 5747 3115 5750
rect 7200 5720 8000 5750
rect 3325 5674 3391 5677
rect 3325 5672 7114 5674
rect 3325 5616 3330 5672
rect 3386 5616 7114 5672
rect 3325 5614 7114 5616
rect 3325 5611 3391 5614
rect 7054 5538 7114 5614
rect 7200 5538 8000 5568
rect 7054 5478 8000 5538
rect 2372 5472 2688 5473
rect 2372 5408 2378 5472
rect 2442 5408 2458 5472
rect 2522 5408 2538 5472
rect 2602 5408 2618 5472
rect 2682 5408 2688 5472
rect 2372 5407 2688 5408
rect 3798 5472 4114 5473
rect 3798 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4114 5472
rect 3798 5407 4114 5408
rect 5224 5472 5540 5473
rect 5224 5408 5230 5472
rect 5294 5408 5310 5472
rect 5374 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5540 5472
rect 5224 5407 5540 5408
rect 6650 5472 6966 5473
rect 6650 5408 6656 5472
rect 6720 5408 6736 5472
rect 6800 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6966 5472
rect 7200 5448 8000 5478
rect 6650 5407 6966 5408
rect 3601 5266 3667 5269
rect 5349 5266 5415 5269
rect 3601 5264 5415 5266
rect 3601 5208 3606 5264
rect 3662 5208 5354 5264
rect 5410 5208 5415 5264
rect 3601 5206 5415 5208
rect 3601 5203 3667 5206
rect 5349 5203 5415 5206
rect 5717 5266 5783 5269
rect 7200 5266 8000 5296
rect 5717 5264 8000 5266
rect 5717 5208 5722 5264
rect 5778 5208 8000 5264
rect 5717 5206 8000 5208
rect 5717 5203 5783 5206
rect 7200 5176 8000 5206
rect 3325 5130 3391 5133
rect 4981 5130 5047 5133
rect 5441 5130 5507 5133
rect 3325 5128 5507 5130
rect 3325 5072 3330 5128
rect 3386 5072 4986 5128
rect 5042 5072 5446 5128
rect 5502 5072 5507 5128
rect 3325 5070 5507 5072
rect 3325 5067 3391 5070
rect 4981 5067 5047 5070
rect 5441 5067 5507 5070
rect 5582 5070 6378 5130
rect 0 4994 800 5024
rect 933 4994 999 4997
rect 0 4992 999 4994
rect 0 4936 938 4992
rect 994 4936 999 4992
rect 0 4934 999 4936
rect 0 4904 800 4934
rect 933 4931 999 4934
rect 5257 4994 5323 4997
rect 5582 4994 5642 5070
rect 5257 4992 5642 4994
rect 5257 4936 5262 4992
rect 5318 4936 5642 4992
rect 5257 4934 5642 4936
rect 6318 4994 6378 5070
rect 7200 4994 8000 5024
rect 6318 4934 8000 4994
rect 5257 4931 5323 4934
rect 1659 4928 1975 4929
rect 1659 4864 1665 4928
rect 1729 4864 1745 4928
rect 1809 4864 1825 4928
rect 1889 4864 1905 4928
rect 1969 4864 1975 4928
rect 1659 4863 1975 4864
rect 3085 4928 3401 4929
rect 3085 4864 3091 4928
rect 3155 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3401 4928
rect 3085 4863 3401 4864
rect 4511 4928 4827 4929
rect 4511 4864 4517 4928
rect 4581 4864 4597 4928
rect 4661 4864 4677 4928
rect 4741 4864 4757 4928
rect 4821 4864 4827 4928
rect 4511 4863 4827 4864
rect 5937 4928 6253 4929
rect 5937 4864 5943 4928
rect 6007 4864 6023 4928
rect 6087 4864 6103 4928
rect 6167 4864 6183 4928
rect 6247 4864 6253 4928
rect 7200 4904 8000 4934
rect 5937 4863 6253 4864
rect 4061 4722 4127 4725
rect 7200 4722 8000 4752
rect 4061 4720 8000 4722
rect 4061 4664 4066 4720
rect 4122 4664 8000 4720
rect 4061 4662 8000 4664
rect 4061 4659 4127 4662
rect 7200 4632 8000 4662
rect 2957 4586 3023 4589
rect 2957 4584 7114 4586
rect 2957 4528 2962 4584
rect 3018 4528 7114 4584
rect 2957 4526 7114 4528
rect 2957 4523 3023 4526
rect 7054 4450 7114 4526
rect 7200 4450 8000 4480
rect 7054 4390 8000 4450
rect 2372 4384 2688 4385
rect 2372 4320 2378 4384
rect 2442 4320 2458 4384
rect 2522 4320 2538 4384
rect 2602 4320 2618 4384
rect 2682 4320 2688 4384
rect 2372 4319 2688 4320
rect 3798 4384 4114 4385
rect 3798 4320 3804 4384
rect 3868 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4114 4384
rect 3798 4319 4114 4320
rect 5224 4384 5540 4385
rect 5224 4320 5230 4384
rect 5294 4320 5310 4384
rect 5374 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5540 4384
rect 5224 4319 5540 4320
rect 6650 4384 6966 4385
rect 6650 4320 6656 4384
rect 6720 4320 6736 4384
rect 6800 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6966 4384
rect 7200 4360 8000 4390
rect 6650 4319 6966 4320
rect 4061 4178 4127 4181
rect 7200 4178 8000 4208
rect 4061 4176 8000 4178
rect 4061 4120 4066 4176
rect 4122 4120 8000 4176
rect 4061 4118 8000 4120
rect 4061 4115 4127 4118
rect 7200 4088 8000 4118
rect 3049 4042 3115 4045
rect 5809 4042 5875 4045
rect 3049 4040 5875 4042
rect 3049 3984 3054 4040
rect 3110 3984 5814 4040
rect 5870 3984 5875 4040
rect 3049 3982 5875 3984
rect 3049 3979 3115 3982
rect 5809 3979 5875 3982
rect 6361 3906 6427 3909
rect 7200 3906 8000 3936
rect 6361 3904 8000 3906
rect 6361 3848 6366 3904
rect 6422 3848 8000 3904
rect 6361 3846 8000 3848
rect 6361 3843 6427 3846
rect 1659 3840 1975 3841
rect 1659 3776 1665 3840
rect 1729 3776 1745 3840
rect 1809 3776 1825 3840
rect 1889 3776 1905 3840
rect 1969 3776 1975 3840
rect 1659 3775 1975 3776
rect 3085 3840 3401 3841
rect 3085 3776 3091 3840
rect 3155 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3401 3840
rect 3085 3775 3401 3776
rect 4511 3840 4827 3841
rect 4511 3776 4517 3840
rect 4581 3776 4597 3840
rect 4661 3776 4677 3840
rect 4741 3776 4757 3840
rect 4821 3776 4827 3840
rect 4511 3775 4827 3776
rect 5937 3840 6253 3841
rect 5937 3776 5943 3840
rect 6007 3776 6023 3840
rect 6087 3776 6103 3840
rect 6167 3776 6183 3840
rect 6247 3776 6253 3840
rect 7200 3816 8000 3846
rect 5937 3775 6253 3776
rect 4061 3634 4127 3637
rect 7200 3634 8000 3664
rect 4061 3632 8000 3634
rect 4061 3576 4066 3632
rect 4122 3576 8000 3632
rect 4061 3574 8000 3576
rect 4061 3571 4127 3574
rect 7200 3544 8000 3574
rect 4061 3498 4127 3501
rect 4061 3496 7114 3498
rect 4061 3440 4066 3496
rect 4122 3440 7114 3496
rect 4061 3438 7114 3440
rect 4061 3435 4127 3438
rect 7054 3362 7114 3438
rect 7200 3362 8000 3392
rect 7054 3302 8000 3362
rect 2372 3296 2688 3297
rect 2372 3232 2378 3296
rect 2442 3232 2458 3296
rect 2522 3232 2538 3296
rect 2602 3232 2618 3296
rect 2682 3232 2688 3296
rect 2372 3231 2688 3232
rect 3798 3296 4114 3297
rect 3798 3232 3804 3296
rect 3868 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4114 3296
rect 3798 3231 4114 3232
rect 5224 3296 5540 3297
rect 5224 3232 5230 3296
rect 5294 3232 5310 3296
rect 5374 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5540 3296
rect 5224 3231 5540 3232
rect 6650 3296 6966 3297
rect 6650 3232 6656 3296
rect 6720 3232 6736 3296
rect 6800 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6966 3296
rect 7200 3272 8000 3302
rect 6650 3231 6966 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 6177 3090 6243 3093
rect 7200 3090 8000 3120
rect 6177 3088 8000 3090
rect 6177 3032 6182 3088
rect 6238 3032 8000 3088
rect 6177 3030 8000 3032
rect 6177 3027 6243 3030
rect 7200 3000 8000 3030
rect 4889 2954 4955 2957
rect 4889 2952 6378 2954
rect 4889 2896 4894 2952
rect 4950 2896 6378 2952
rect 4889 2894 6378 2896
rect 4889 2891 4955 2894
rect 6318 2818 6378 2894
rect 7200 2818 8000 2848
rect 6318 2758 8000 2818
rect 1659 2752 1975 2753
rect 1659 2688 1665 2752
rect 1729 2688 1745 2752
rect 1809 2688 1825 2752
rect 1889 2688 1905 2752
rect 1969 2688 1975 2752
rect 1659 2687 1975 2688
rect 3085 2752 3401 2753
rect 3085 2688 3091 2752
rect 3155 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3401 2752
rect 3085 2687 3401 2688
rect 4511 2752 4827 2753
rect 4511 2688 4517 2752
rect 4581 2688 4597 2752
rect 4661 2688 4677 2752
rect 4741 2688 4757 2752
rect 4821 2688 4827 2752
rect 4511 2687 4827 2688
rect 5937 2752 6253 2753
rect 5937 2688 5943 2752
rect 6007 2688 6023 2752
rect 6087 2688 6103 2752
rect 6167 2688 6183 2752
rect 6247 2688 6253 2752
rect 7200 2728 8000 2758
rect 5937 2687 6253 2688
rect 4429 2546 4495 2549
rect 7200 2546 8000 2576
rect 4429 2544 8000 2546
rect 4429 2488 4434 2544
rect 4490 2488 8000 2544
rect 4429 2486 8000 2488
rect 4429 2483 4495 2486
rect 7200 2456 8000 2486
rect 6177 2410 6243 2413
rect 6177 2408 7114 2410
rect 6177 2352 6182 2408
rect 6238 2352 7114 2408
rect 6177 2350 7114 2352
rect 6177 2347 6243 2350
rect 7054 2274 7114 2350
rect 7200 2274 8000 2304
rect 7054 2214 8000 2274
rect 2372 2208 2688 2209
rect 2372 2144 2378 2208
rect 2442 2144 2458 2208
rect 2522 2144 2538 2208
rect 2602 2144 2618 2208
rect 2682 2144 2688 2208
rect 2372 2143 2688 2144
rect 3798 2208 4114 2209
rect 3798 2144 3804 2208
rect 3868 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4114 2208
rect 3798 2143 4114 2144
rect 5224 2208 5540 2209
rect 5224 2144 5230 2208
rect 5294 2144 5310 2208
rect 5374 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5540 2208
rect 5224 2143 5540 2144
rect 6650 2208 6966 2209
rect 6650 2144 6656 2208
rect 6720 2144 6736 2208
rect 6800 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6966 2208
rect 7200 2184 8000 2214
rect 6650 2143 6966 2144
rect 1577 2038 1643 2041
rect 798 2036 1643 2038
rect 798 1980 1582 2036
rect 1638 1980 1643 2036
rect 798 1978 1643 1980
rect 798 1932 858 1978
rect 1577 1975 1643 1978
rect 0 1842 858 1932
rect 7200 1912 8000 2032
rect 0 1812 800 1842
<< via3 >>
rect 2378 5468 2442 5472
rect 2378 5412 2382 5468
rect 2382 5412 2438 5468
rect 2438 5412 2442 5468
rect 2378 5408 2442 5412
rect 2458 5468 2522 5472
rect 2458 5412 2462 5468
rect 2462 5412 2518 5468
rect 2518 5412 2522 5468
rect 2458 5408 2522 5412
rect 2538 5468 2602 5472
rect 2538 5412 2542 5468
rect 2542 5412 2598 5468
rect 2598 5412 2602 5468
rect 2538 5408 2602 5412
rect 2618 5468 2682 5472
rect 2618 5412 2622 5468
rect 2622 5412 2678 5468
rect 2678 5412 2682 5468
rect 2618 5408 2682 5412
rect 3804 5468 3868 5472
rect 3804 5412 3808 5468
rect 3808 5412 3864 5468
rect 3864 5412 3868 5468
rect 3804 5408 3868 5412
rect 3884 5468 3948 5472
rect 3884 5412 3888 5468
rect 3888 5412 3944 5468
rect 3944 5412 3948 5468
rect 3884 5408 3948 5412
rect 3964 5468 4028 5472
rect 3964 5412 3968 5468
rect 3968 5412 4024 5468
rect 4024 5412 4028 5468
rect 3964 5408 4028 5412
rect 4044 5468 4108 5472
rect 4044 5412 4048 5468
rect 4048 5412 4104 5468
rect 4104 5412 4108 5468
rect 4044 5408 4108 5412
rect 5230 5468 5294 5472
rect 5230 5412 5234 5468
rect 5234 5412 5290 5468
rect 5290 5412 5294 5468
rect 5230 5408 5294 5412
rect 5310 5468 5374 5472
rect 5310 5412 5314 5468
rect 5314 5412 5370 5468
rect 5370 5412 5374 5468
rect 5310 5408 5374 5412
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 6656 5468 6720 5472
rect 6656 5412 6660 5468
rect 6660 5412 6716 5468
rect 6716 5412 6720 5468
rect 6656 5408 6720 5412
rect 6736 5468 6800 5472
rect 6736 5412 6740 5468
rect 6740 5412 6796 5468
rect 6796 5412 6800 5468
rect 6736 5408 6800 5412
rect 6816 5468 6880 5472
rect 6816 5412 6820 5468
rect 6820 5412 6876 5468
rect 6876 5412 6880 5468
rect 6816 5408 6880 5412
rect 6896 5468 6960 5472
rect 6896 5412 6900 5468
rect 6900 5412 6956 5468
rect 6956 5412 6960 5468
rect 6896 5408 6960 5412
rect 1665 4924 1729 4928
rect 1665 4868 1669 4924
rect 1669 4868 1725 4924
rect 1725 4868 1729 4924
rect 1665 4864 1729 4868
rect 1745 4924 1809 4928
rect 1745 4868 1749 4924
rect 1749 4868 1805 4924
rect 1805 4868 1809 4924
rect 1745 4864 1809 4868
rect 1825 4924 1889 4928
rect 1825 4868 1829 4924
rect 1829 4868 1885 4924
rect 1885 4868 1889 4924
rect 1825 4864 1889 4868
rect 1905 4924 1969 4928
rect 1905 4868 1909 4924
rect 1909 4868 1965 4924
rect 1965 4868 1969 4924
rect 1905 4864 1969 4868
rect 3091 4924 3155 4928
rect 3091 4868 3095 4924
rect 3095 4868 3151 4924
rect 3151 4868 3155 4924
rect 3091 4864 3155 4868
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 4517 4924 4581 4928
rect 4517 4868 4521 4924
rect 4521 4868 4577 4924
rect 4577 4868 4581 4924
rect 4517 4864 4581 4868
rect 4597 4924 4661 4928
rect 4597 4868 4601 4924
rect 4601 4868 4657 4924
rect 4657 4868 4661 4924
rect 4597 4864 4661 4868
rect 4677 4924 4741 4928
rect 4677 4868 4681 4924
rect 4681 4868 4737 4924
rect 4737 4868 4741 4924
rect 4677 4864 4741 4868
rect 4757 4924 4821 4928
rect 4757 4868 4761 4924
rect 4761 4868 4817 4924
rect 4817 4868 4821 4924
rect 4757 4864 4821 4868
rect 5943 4924 6007 4928
rect 5943 4868 5947 4924
rect 5947 4868 6003 4924
rect 6003 4868 6007 4924
rect 5943 4864 6007 4868
rect 6023 4924 6087 4928
rect 6023 4868 6027 4924
rect 6027 4868 6083 4924
rect 6083 4868 6087 4924
rect 6023 4864 6087 4868
rect 6103 4924 6167 4928
rect 6103 4868 6107 4924
rect 6107 4868 6163 4924
rect 6163 4868 6167 4924
rect 6103 4864 6167 4868
rect 6183 4924 6247 4928
rect 6183 4868 6187 4924
rect 6187 4868 6243 4924
rect 6243 4868 6247 4924
rect 6183 4864 6247 4868
rect 2378 4380 2442 4384
rect 2378 4324 2382 4380
rect 2382 4324 2438 4380
rect 2438 4324 2442 4380
rect 2378 4320 2442 4324
rect 2458 4380 2522 4384
rect 2458 4324 2462 4380
rect 2462 4324 2518 4380
rect 2518 4324 2522 4380
rect 2458 4320 2522 4324
rect 2538 4380 2602 4384
rect 2538 4324 2542 4380
rect 2542 4324 2598 4380
rect 2598 4324 2602 4380
rect 2538 4320 2602 4324
rect 2618 4380 2682 4384
rect 2618 4324 2622 4380
rect 2622 4324 2678 4380
rect 2678 4324 2682 4380
rect 2618 4320 2682 4324
rect 3804 4380 3868 4384
rect 3804 4324 3808 4380
rect 3808 4324 3864 4380
rect 3864 4324 3868 4380
rect 3804 4320 3868 4324
rect 3884 4380 3948 4384
rect 3884 4324 3888 4380
rect 3888 4324 3944 4380
rect 3944 4324 3948 4380
rect 3884 4320 3948 4324
rect 3964 4380 4028 4384
rect 3964 4324 3968 4380
rect 3968 4324 4024 4380
rect 4024 4324 4028 4380
rect 3964 4320 4028 4324
rect 4044 4380 4108 4384
rect 4044 4324 4048 4380
rect 4048 4324 4104 4380
rect 4104 4324 4108 4380
rect 4044 4320 4108 4324
rect 5230 4380 5294 4384
rect 5230 4324 5234 4380
rect 5234 4324 5290 4380
rect 5290 4324 5294 4380
rect 5230 4320 5294 4324
rect 5310 4380 5374 4384
rect 5310 4324 5314 4380
rect 5314 4324 5370 4380
rect 5370 4324 5374 4380
rect 5310 4320 5374 4324
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 6656 4380 6720 4384
rect 6656 4324 6660 4380
rect 6660 4324 6716 4380
rect 6716 4324 6720 4380
rect 6656 4320 6720 4324
rect 6736 4380 6800 4384
rect 6736 4324 6740 4380
rect 6740 4324 6796 4380
rect 6796 4324 6800 4380
rect 6736 4320 6800 4324
rect 6816 4380 6880 4384
rect 6816 4324 6820 4380
rect 6820 4324 6876 4380
rect 6876 4324 6880 4380
rect 6816 4320 6880 4324
rect 6896 4380 6960 4384
rect 6896 4324 6900 4380
rect 6900 4324 6956 4380
rect 6956 4324 6960 4380
rect 6896 4320 6960 4324
rect 1665 3836 1729 3840
rect 1665 3780 1669 3836
rect 1669 3780 1725 3836
rect 1725 3780 1729 3836
rect 1665 3776 1729 3780
rect 1745 3836 1809 3840
rect 1745 3780 1749 3836
rect 1749 3780 1805 3836
rect 1805 3780 1809 3836
rect 1745 3776 1809 3780
rect 1825 3836 1889 3840
rect 1825 3780 1829 3836
rect 1829 3780 1885 3836
rect 1885 3780 1889 3836
rect 1825 3776 1889 3780
rect 1905 3836 1969 3840
rect 1905 3780 1909 3836
rect 1909 3780 1965 3836
rect 1965 3780 1969 3836
rect 1905 3776 1969 3780
rect 3091 3836 3155 3840
rect 3091 3780 3095 3836
rect 3095 3780 3151 3836
rect 3151 3780 3155 3836
rect 3091 3776 3155 3780
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 4517 3836 4581 3840
rect 4517 3780 4521 3836
rect 4521 3780 4577 3836
rect 4577 3780 4581 3836
rect 4517 3776 4581 3780
rect 4597 3836 4661 3840
rect 4597 3780 4601 3836
rect 4601 3780 4657 3836
rect 4657 3780 4661 3836
rect 4597 3776 4661 3780
rect 4677 3836 4741 3840
rect 4677 3780 4681 3836
rect 4681 3780 4737 3836
rect 4737 3780 4741 3836
rect 4677 3776 4741 3780
rect 4757 3836 4821 3840
rect 4757 3780 4761 3836
rect 4761 3780 4817 3836
rect 4817 3780 4821 3836
rect 4757 3776 4821 3780
rect 5943 3836 6007 3840
rect 5943 3780 5947 3836
rect 5947 3780 6003 3836
rect 6003 3780 6007 3836
rect 5943 3776 6007 3780
rect 6023 3836 6087 3840
rect 6023 3780 6027 3836
rect 6027 3780 6083 3836
rect 6083 3780 6087 3836
rect 6023 3776 6087 3780
rect 6103 3836 6167 3840
rect 6103 3780 6107 3836
rect 6107 3780 6163 3836
rect 6163 3780 6167 3836
rect 6103 3776 6167 3780
rect 6183 3836 6247 3840
rect 6183 3780 6187 3836
rect 6187 3780 6243 3836
rect 6243 3780 6247 3836
rect 6183 3776 6247 3780
rect 2378 3292 2442 3296
rect 2378 3236 2382 3292
rect 2382 3236 2438 3292
rect 2438 3236 2442 3292
rect 2378 3232 2442 3236
rect 2458 3292 2522 3296
rect 2458 3236 2462 3292
rect 2462 3236 2518 3292
rect 2518 3236 2522 3292
rect 2458 3232 2522 3236
rect 2538 3292 2602 3296
rect 2538 3236 2542 3292
rect 2542 3236 2598 3292
rect 2598 3236 2602 3292
rect 2538 3232 2602 3236
rect 2618 3292 2682 3296
rect 2618 3236 2622 3292
rect 2622 3236 2678 3292
rect 2678 3236 2682 3292
rect 2618 3232 2682 3236
rect 3804 3292 3868 3296
rect 3804 3236 3808 3292
rect 3808 3236 3864 3292
rect 3864 3236 3868 3292
rect 3804 3232 3868 3236
rect 3884 3292 3948 3296
rect 3884 3236 3888 3292
rect 3888 3236 3944 3292
rect 3944 3236 3948 3292
rect 3884 3232 3948 3236
rect 3964 3292 4028 3296
rect 3964 3236 3968 3292
rect 3968 3236 4024 3292
rect 4024 3236 4028 3292
rect 3964 3232 4028 3236
rect 4044 3292 4108 3296
rect 4044 3236 4048 3292
rect 4048 3236 4104 3292
rect 4104 3236 4108 3292
rect 4044 3232 4108 3236
rect 5230 3292 5294 3296
rect 5230 3236 5234 3292
rect 5234 3236 5290 3292
rect 5290 3236 5294 3292
rect 5230 3232 5294 3236
rect 5310 3292 5374 3296
rect 5310 3236 5314 3292
rect 5314 3236 5370 3292
rect 5370 3236 5374 3292
rect 5310 3232 5374 3236
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 6656 3292 6720 3296
rect 6656 3236 6660 3292
rect 6660 3236 6716 3292
rect 6716 3236 6720 3292
rect 6656 3232 6720 3236
rect 6736 3292 6800 3296
rect 6736 3236 6740 3292
rect 6740 3236 6796 3292
rect 6796 3236 6800 3292
rect 6736 3232 6800 3236
rect 6816 3292 6880 3296
rect 6816 3236 6820 3292
rect 6820 3236 6876 3292
rect 6876 3236 6880 3292
rect 6816 3232 6880 3236
rect 6896 3292 6960 3296
rect 6896 3236 6900 3292
rect 6900 3236 6956 3292
rect 6956 3236 6960 3292
rect 6896 3232 6960 3236
rect 1665 2748 1729 2752
rect 1665 2692 1669 2748
rect 1669 2692 1725 2748
rect 1725 2692 1729 2748
rect 1665 2688 1729 2692
rect 1745 2748 1809 2752
rect 1745 2692 1749 2748
rect 1749 2692 1805 2748
rect 1805 2692 1809 2748
rect 1745 2688 1809 2692
rect 1825 2748 1889 2752
rect 1825 2692 1829 2748
rect 1829 2692 1885 2748
rect 1885 2692 1889 2748
rect 1825 2688 1889 2692
rect 1905 2748 1969 2752
rect 1905 2692 1909 2748
rect 1909 2692 1965 2748
rect 1965 2692 1969 2748
rect 1905 2688 1969 2692
rect 3091 2748 3155 2752
rect 3091 2692 3095 2748
rect 3095 2692 3151 2748
rect 3151 2692 3155 2748
rect 3091 2688 3155 2692
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 4517 2748 4581 2752
rect 4517 2692 4521 2748
rect 4521 2692 4577 2748
rect 4577 2692 4581 2748
rect 4517 2688 4581 2692
rect 4597 2748 4661 2752
rect 4597 2692 4601 2748
rect 4601 2692 4657 2748
rect 4657 2692 4661 2748
rect 4597 2688 4661 2692
rect 4677 2748 4741 2752
rect 4677 2692 4681 2748
rect 4681 2692 4737 2748
rect 4737 2692 4741 2748
rect 4677 2688 4741 2692
rect 4757 2748 4821 2752
rect 4757 2692 4761 2748
rect 4761 2692 4817 2748
rect 4817 2692 4821 2748
rect 4757 2688 4821 2692
rect 5943 2748 6007 2752
rect 5943 2692 5947 2748
rect 5947 2692 6003 2748
rect 6003 2692 6007 2748
rect 5943 2688 6007 2692
rect 6023 2748 6087 2752
rect 6023 2692 6027 2748
rect 6027 2692 6083 2748
rect 6083 2692 6087 2748
rect 6023 2688 6087 2692
rect 6103 2748 6167 2752
rect 6103 2692 6107 2748
rect 6107 2692 6163 2748
rect 6163 2692 6167 2748
rect 6103 2688 6167 2692
rect 6183 2748 6247 2752
rect 6183 2692 6187 2748
rect 6187 2692 6243 2748
rect 6243 2692 6247 2748
rect 6183 2688 6247 2692
rect 2378 2204 2442 2208
rect 2378 2148 2382 2204
rect 2382 2148 2438 2204
rect 2438 2148 2442 2204
rect 2378 2144 2442 2148
rect 2458 2204 2522 2208
rect 2458 2148 2462 2204
rect 2462 2148 2518 2204
rect 2518 2148 2522 2204
rect 2458 2144 2522 2148
rect 2538 2204 2602 2208
rect 2538 2148 2542 2204
rect 2542 2148 2598 2204
rect 2598 2148 2602 2204
rect 2538 2144 2602 2148
rect 2618 2204 2682 2208
rect 2618 2148 2622 2204
rect 2622 2148 2678 2204
rect 2678 2148 2682 2204
rect 2618 2144 2682 2148
rect 3804 2204 3868 2208
rect 3804 2148 3808 2204
rect 3808 2148 3864 2204
rect 3864 2148 3868 2204
rect 3804 2144 3868 2148
rect 3884 2204 3948 2208
rect 3884 2148 3888 2204
rect 3888 2148 3944 2204
rect 3944 2148 3948 2204
rect 3884 2144 3948 2148
rect 3964 2204 4028 2208
rect 3964 2148 3968 2204
rect 3968 2148 4024 2204
rect 4024 2148 4028 2204
rect 3964 2144 4028 2148
rect 4044 2204 4108 2208
rect 4044 2148 4048 2204
rect 4048 2148 4104 2204
rect 4104 2148 4108 2204
rect 4044 2144 4108 2148
rect 5230 2204 5294 2208
rect 5230 2148 5234 2204
rect 5234 2148 5290 2204
rect 5290 2148 5294 2204
rect 5230 2144 5294 2148
rect 5310 2204 5374 2208
rect 5310 2148 5314 2204
rect 5314 2148 5370 2204
rect 5370 2148 5374 2204
rect 5310 2144 5374 2148
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 6656 2204 6720 2208
rect 6656 2148 6660 2204
rect 6660 2148 6716 2204
rect 6716 2148 6720 2204
rect 6656 2144 6720 2148
rect 6736 2204 6800 2208
rect 6736 2148 6740 2204
rect 6740 2148 6796 2204
rect 6796 2148 6800 2204
rect 6736 2144 6800 2148
rect 6816 2204 6880 2208
rect 6816 2148 6820 2204
rect 6820 2148 6876 2204
rect 6876 2148 6880 2204
rect 6816 2144 6880 2148
rect 6896 2204 6960 2208
rect 6896 2148 6900 2204
rect 6900 2148 6956 2204
rect 6956 2148 6960 2204
rect 6896 2144 6960 2148
<< metal4 >>
rect 1657 4928 1977 5488
rect 1657 4864 1665 4928
rect 1729 4864 1745 4928
rect 1809 4864 1825 4928
rect 1889 4864 1905 4928
rect 1969 4864 1977 4928
rect 1657 3840 1977 4864
rect 1657 3776 1665 3840
rect 1729 3776 1745 3840
rect 1809 3776 1825 3840
rect 1889 3776 1905 3840
rect 1969 3776 1977 3840
rect 1657 2752 1977 3776
rect 1657 2688 1665 2752
rect 1729 2688 1745 2752
rect 1809 2688 1825 2752
rect 1889 2688 1905 2752
rect 1969 2688 1977 2752
rect 1657 2128 1977 2688
rect 2370 5472 2690 5488
rect 2370 5408 2378 5472
rect 2442 5408 2458 5472
rect 2522 5408 2538 5472
rect 2602 5408 2618 5472
rect 2682 5408 2690 5472
rect 2370 4384 2690 5408
rect 2370 4320 2378 4384
rect 2442 4320 2458 4384
rect 2522 4320 2538 4384
rect 2602 4320 2618 4384
rect 2682 4320 2690 4384
rect 2370 3296 2690 4320
rect 2370 3232 2378 3296
rect 2442 3232 2458 3296
rect 2522 3232 2538 3296
rect 2602 3232 2618 3296
rect 2682 3232 2690 3296
rect 2370 2208 2690 3232
rect 2370 2144 2378 2208
rect 2442 2144 2458 2208
rect 2522 2144 2538 2208
rect 2602 2144 2618 2208
rect 2682 2144 2690 2208
rect 2370 2128 2690 2144
rect 3083 4928 3403 5488
rect 3083 4864 3091 4928
rect 3155 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3403 4928
rect 3083 3840 3403 4864
rect 3083 3776 3091 3840
rect 3155 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3403 3840
rect 3083 2752 3403 3776
rect 3083 2688 3091 2752
rect 3155 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3403 2752
rect 3083 2128 3403 2688
rect 3796 5472 4116 5488
rect 3796 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4116 5472
rect 3796 4384 4116 5408
rect 3796 4320 3804 4384
rect 3868 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4116 4384
rect 3796 3296 4116 4320
rect 3796 3232 3804 3296
rect 3868 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4116 3296
rect 3796 2208 4116 3232
rect 3796 2144 3804 2208
rect 3868 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4116 2208
rect 3796 2128 4116 2144
rect 4509 4928 4829 5488
rect 4509 4864 4517 4928
rect 4581 4864 4597 4928
rect 4661 4864 4677 4928
rect 4741 4864 4757 4928
rect 4821 4864 4829 4928
rect 4509 3840 4829 4864
rect 4509 3776 4517 3840
rect 4581 3776 4597 3840
rect 4661 3776 4677 3840
rect 4741 3776 4757 3840
rect 4821 3776 4829 3840
rect 4509 2752 4829 3776
rect 4509 2688 4517 2752
rect 4581 2688 4597 2752
rect 4661 2688 4677 2752
rect 4741 2688 4757 2752
rect 4821 2688 4829 2752
rect 4509 2128 4829 2688
rect 5222 5472 5542 5488
rect 5222 5408 5230 5472
rect 5294 5408 5310 5472
rect 5374 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5542 5472
rect 5222 4384 5542 5408
rect 5222 4320 5230 4384
rect 5294 4320 5310 4384
rect 5374 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5542 4384
rect 5222 3296 5542 4320
rect 5222 3232 5230 3296
rect 5294 3232 5310 3296
rect 5374 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5542 3296
rect 5222 2208 5542 3232
rect 5222 2144 5230 2208
rect 5294 2144 5310 2208
rect 5374 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5542 2208
rect 5222 2128 5542 2144
rect 5935 4928 6255 5488
rect 5935 4864 5943 4928
rect 6007 4864 6023 4928
rect 6087 4864 6103 4928
rect 6167 4864 6183 4928
rect 6247 4864 6255 4928
rect 5935 3840 6255 4864
rect 5935 3776 5943 3840
rect 6007 3776 6023 3840
rect 6087 3776 6103 3840
rect 6167 3776 6183 3840
rect 6247 3776 6255 3840
rect 5935 2752 6255 3776
rect 5935 2688 5943 2752
rect 6007 2688 6023 2752
rect 6087 2688 6103 2752
rect 6167 2688 6183 2752
rect 6247 2688 6255 2752
rect 5935 2128 6255 2688
rect 6648 5472 6968 5488
rect 6648 5408 6656 5472
rect 6720 5408 6736 5472
rect 6800 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6968 5472
rect 6648 4384 6968 5408
rect 6648 4320 6656 4384
rect 6720 4320 6736 4384
rect 6800 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6968 4384
rect 6648 3296 6968 4320
rect 6648 3232 6656 3296
rect 6720 3232 6736 3296
rect 6800 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6968 3296
rect 6648 2208 6968 3232
rect 6648 2144 6656 2208
rect 6720 2144 6736 2208
rect 6800 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6968 2208
rect 6648 2128 6968 2144
use sky130_fd_sc_hd__inv_2  _16_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _17_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform -1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _18_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _19_
timestamp 1733649010
transform -1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _20_
timestamp 1733649010
transform -1 0 5980 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _21_
timestamp 1733649010
transform 1 0 5520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _22_
timestamp 1733649010
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _23_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _24_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _25_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform -1 0 6072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 1733649010
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _27_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 4600 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _28_
timestamp 1733649010
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _29_
timestamp 1733649010
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _30_
timestamp 1733649010
transform 1 0 4140 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _31_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform -1 0 4416 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _32_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 5428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _33_
timestamp 1733649010
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _34_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 4784 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _35_ ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 4784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1733649010
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_37 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1733649010
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1733649010
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1733649010
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_33
timestamp 1733649010
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1733649010
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1733649010
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1733649010
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1733649010
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1733649010
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1733649010
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 1733649010
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_44
timestamp 1733649010
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1733649010
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_38
timestamp 1733649010
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_29
timestamp 1733649010
transform 1 0 3772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1733649010
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1733649010
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1733649010
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1733649010
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1733649010
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1733649010
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1733649010
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1733649010
transform -1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1733649010
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1733649010
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1733649010
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1733649010
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1733649010
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1733649010
transform -1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output16 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform -1 0 2852 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output17
timestamp 1733649010
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output18
timestamp 1733649010
transform -1 0 2852 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output19
timestamp 1733649010
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1733649010
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1733649010
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1733649010
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1733649010
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1733649010
transform -1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1733649010
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1733649010
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1733649010
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1733649010
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1733649010
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1733649010
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold
timestamp 1733649010
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1733649010
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1733649010
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1733649010
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1733649010
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1733649010
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1733649010
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1733649010
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
<< labels >>
flabel metal4 s 6648 2128 6968 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5222 2128 5542 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3796 2128 4116 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2370 2128 2690 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5935 2128 6255 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4509 2128 4829 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3083 2128 3403 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1657 2128 1977 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 7200 1912 8000 2032 0 FreeSans 600 0 0 0 in0
port 3 nsew
flabel metal3 s 7200 2184 8000 2304 0 FreeSans 600 0 0 0 in1
port 4 nsew
flabel metal3 s 7200 4632 8000 4752 0 FreeSans 600 0 0 0 in10
port 5 nsew
flabel metal3 s 7200 4904 8000 5024 0 FreeSans 600 0 0 0 in11
port 6 nsew
flabel metal3 s 7200 5176 8000 5296 0 FreeSans 600 0 0 0 in12
port 7 nsew
flabel metal3 s 7200 5448 8000 5568 0 FreeSans 600 0 0 0 in13
port 8 nsew
flabel metal3 s 7200 5720 8000 5840 0 FreeSans 600 0 0 0 in14
port 9 nsew
flabel metal3 s 7200 5992 8000 6112 0 FreeSans 600 0 0 0 in15
port 10 nsew
flabel metal3 s 7200 2456 8000 2576 0 FreeSans 600 0 0 0 in2
port 11 nsew
flabel metal3 s 7200 2728 8000 2848 0 FreeSans 600 0 0 0 in3
port 12 nsew
flabel metal3 s 7200 3000 8000 3120 0 FreeSans 600 0 0 0 in4
port 13 nsew
flabel metal3 s 7200 3272 8000 3392 0 FreeSans 600 0 0 0 in5
port 14 nsew
flabel metal3 s 7200 3544 8000 3664 0 FreeSans 600 0 0 0 in6
port 15 nsew
flabel metal3 s 7200 3816 8000 3936 0 FreeSans 600 0 0 0 in7
port 16 nsew
flabel metal3 s 7200 4088 8000 4208 0 FreeSans 600 0 0 0 in8
port 17 nsew
flabel metal3 s 7200 4360 8000 4480 0 FreeSans 600 0 0 0 in9
port 18 nsew
flabel metal3 s 0 3000 800 3120 0 FreeSans 600 0 0 0 out[1]
port 20 nsew
flabel metal3 s 0 4904 800 5024 0 FreeSans 600 0 0 0 out[2]
port 21 nsew
flabel metal3 s 0 5720 800 5840 0 FreeSans 600 0 0 0 out[3]
port 22 nsew
flabel metal3 s 0 1812 800 1932 0 FreeSans 600 0 0 0 out[0]
port 19 nsew
<< properties >>
string FIXED_BBOX 0 0 8000 8000
<< end >>
