magic
tech sky130B
magscale 1 2
timestamp 1732044439
<< error_s >>
rect 251 -6359 309 -6353
rect 531 -6359 589 -6353
rect 811 -6359 869 -6353
rect 1091 -6359 1149 -6353
rect 1371 -6359 1429 -6353
rect 1651 -6359 1709 -6353
rect 1931 -6359 1989 -6353
rect 2211 -6359 2269 -6353
rect 2491 -6359 2549 -6353
rect 2771 -6359 2829 -6353
rect 251 -6393 263 -6359
rect 531 -6393 543 -6359
rect 811 -6393 823 -6359
rect 1091 -6393 1103 -6359
rect 1371 -6393 1383 -6359
rect 1651 -6393 1663 -6359
rect 1931 -6393 1943 -6359
rect 2211 -6393 2223 -6359
rect 2491 -6393 2503 -6359
rect 2771 -6393 2783 -6359
rect 251 -6399 309 -6393
rect 531 -6399 589 -6393
rect 811 -6399 869 -6393
rect 1091 -6399 1149 -6393
rect 1371 -6399 1429 -6393
rect 1651 -6399 1709 -6393
rect 1931 -6399 1989 -6393
rect 2211 -6399 2269 -6393
rect 2491 -6399 2549 -6393
rect 2771 -6399 2829 -6393
rect 598 -7084 618 -7056
rect 626 -7094 646 -7084
rect 670 -7094 690 -7056
rect 251 -7567 309 -7561
rect 531 -7567 589 -7561
rect 811 -7567 869 -7561
rect 1091 -7567 1149 -7561
rect 1371 -7567 1429 -7561
rect 1651 -7567 1709 -7561
rect 1931 -7567 1989 -7561
rect 2211 -7567 2269 -7561
rect 2491 -7567 2549 -7561
rect 2771 -7567 2829 -7561
rect 251 -7601 263 -7567
rect 531 -7601 543 -7567
rect 811 -7601 823 -7567
rect 1091 -7601 1103 -7567
rect 1371 -7601 1383 -7567
rect 1651 -7601 1663 -7567
rect 1931 -7601 1943 -7567
rect 2211 -7601 2223 -7567
rect 2491 -7601 2503 -7567
rect 2771 -7601 2783 -7567
rect 251 -7607 309 -7601
rect 531 -7607 589 -7601
rect 811 -7607 869 -7601
rect 1091 -7607 1149 -7601
rect 1371 -7607 1429 -7601
rect 1651 -7607 1709 -7601
rect 1931 -7607 1989 -7601
rect 2211 -7607 2269 -7601
rect 2491 -7607 2549 -7601
rect 2771 -7607 2829 -7601
<< metal1 >>
rect 254 -6242 306 -6232
rect 254 -6304 306 -6294
rect 534 -6242 586 -6232
rect 534 -6304 586 -6294
rect 1374 -6242 1426 -6232
rect 1374 -6304 1426 -6294
rect 1654 -6242 1706 -6232
rect 1654 -6304 1706 -6294
rect 2494 -6242 2546 -6232
rect 2494 -6304 2546 -6294
rect 2774 -6242 2826 -6232
rect 2774 -6304 2826 -6294
rect 944 -6402 954 -6348
rect 1006 -6402 1016 -6348
rect 2064 -6402 2074 -6348
rect 2126 -6402 2136 -6348
rect 346 -6866 382 -6600
rect 626 -6866 662 -6600
rect 1466 -6866 1502 -6600
rect 1746 -6866 1782 -6600
rect 2586 -6866 2622 -6600
rect 2866 -6866 2902 -6600
rect 338 -6876 390 -6866
rect 338 -6938 390 -6928
rect 618 -6876 670 -6866
rect 618 -6938 670 -6928
rect 1458 -6876 1510 -6866
rect 1458 -6938 1510 -6928
rect 1738 -6876 1790 -6866
rect 1738 -6938 1790 -6928
rect 2578 -6876 2630 -6866
rect 2578 -6938 2630 -6928
rect 2858 -6876 2910 -6866
rect 2858 -6938 2910 -6928
rect 338 -7032 390 -7022
rect 338 -7094 390 -7084
rect 618 -7032 670 -7022
rect 618 -7094 626 -7084
rect 662 -7094 670 -7084
rect 1458 -7032 1510 -7022
rect 1458 -7094 1510 -7084
rect 1738 -7032 1790 -7022
rect 1738 -7094 1790 -7084
rect 2578 -7032 2630 -7022
rect 2578 -7094 2630 -7084
rect 2858 -7032 2910 -7022
rect 2858 -7094 2910 -7084
rect 346 -7360 382 -7094
rect 1466 -7360 1502 -7094
rect 1746 -7360 1782 -7094
rect 2586 -7360 2622 -7094
rect 2866 -7360 2902 -7094
rect 384 -7610 394 -7556
rect 446 -7610 456 -7556
rect 1504 -7610 1514 -7556
rect 1566 -7610 1576 -7556
rect 2624 -7610 2634 -7556
rect 2686 -7610 2696 -7556
rect 814 -7666 866 -7656
rect 814 -7728 866 -7718
rect 1094 -7666 1146 -7656
rect 1094 -7728 1146 -7718
rect 1934 -7666 1986 -7656
rect 1934 -7728 1986 -7718
rect 2214 -7666 2266 -7656
rect 2214 -7728 2266 -7718
<< via1 >>
rect 254 -6294 306 -6242
rect 534 -6294 586 -6242
rect 1374 -6294 1426 -6242
rect 1654 -6294 1706 -6242
rect 2494 -6294 2546 -6242
rect 2774 -6294 2826 -6242
rect 954 -6402 1006 -6348
rect 2074 -6402 2126 -6348
rect 338 -6928 390 -6876
rect 618 -6928 670 -6876
rect 1458 -6928 1510 -6876
rect 1738 -6928 1790 -6876
rect 2578 -6928 2630 -6876
rect 2858 -6928 2910 -6876
rect 338 -7084 390 -7032
rect 618 -7084 670 -7032
rect 1458 -7084 1510 -7032
rect 1738 -7084 1790 -7032
rect 2578 -7084 2630 -7032
rect 2858 -7084 2910 -7032
rect 394 -7610 446 -7556
rect 1514 -7610 1566 -7556
rect 2634 -7610 2686 -7556
rect 814 -7718 866 -7666
rect 1094 -7718 1146 -7666
rect 1934 -7718 1986 -7666
rect 2214 -7718 2266 -7666
<< metal2 >>
rect 244 -6294 254 -6242
rect 306 -6294 316 -6242
rect 524 -6294 534 -6242
rect 586 -6294 596 -6242
rect 1364 -6294 1374 -6242
rect 1426 -6294 1436 -6242
rect 1644 -6294 1654 -6242
rect 1706 -6294 1716 -6242
rect 2484 -6294 2494 -6242
rect 2546 -6294 2556 -6242
rect 2764 -6294 2774 -6242
rect 2826 -6294 2836 -6242
rect 954 -6348 1006 -6338
rect 954 -6412 1006 -6402
rect 2074 -6348 2126 -6338
rect 2074 -6412 2126 -6402
rect 328 -6928 338 -6876
rect 390 -6928 400 -6876
rect 608 -6928 618 -6876
rect 670 -6928 680 -6876
rect 1448 -6928 1458 -6876
rect 1510 -6928 1520 -6876
rect 1728 -6928 1738 -6876
rect 1790 -6928 1800 -6876
rect 2568 -6928 2578 -6876
rect 2630 -6928 2640 -6876
rect 2848 -6928 2858 -6876
rect 2910 -6928 2920 -6876
rect 328 -7084 338 -7032
rect 390 -7084 400 -7032
rect 608 -7084 618 -7032
rect 670 -7084 680 -7032
rect 1448 -7084 1458 -7032
rect 1510 -7084 1520 -7032
rect 1728 -7084 1738 -7032
rect 1790 -7084 1800 -7032
rect 2568 -7084 2578 -7032
rect 2630 -7084 2640 -7032
rect 2848 -7084 2858 -7032
rect 2910 -7084 2920 -7032
rect 394 -7556 446 -7546
rect 394 -7620 446 -7610
rect 1514 -7556 1566 -7546
rect 1514 -7620 1566 -7610
rect 2634 -7556 2686 -7546
rect 2634 -7620 2686 -7610
rect 804 -7718 814 -7666
rect 866 -7718 876 -7666
rect 1084 -7718 1094 -7666
rect 1146 -7718 1156 -7666
rect 1924 -7718 1934 -7666
rect 1986 -7718 1996 -7666
rect 2204 -7718 2214 -7666
rect 2266 -7718 2276 -7666
use sky130_fd_pr__nfet_01v8_72KZQ8  xm49
timestamp 1732044439
transform 1 0 280 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm50
timestamp 1732044439
transform 1 0 560 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm51
timestamp 1732044439
transform 1 0 840 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm52
timestamp 1732044439
transform 1 0 1120 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm53
timestamp 1732044439
transform 1 0 1400 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm54
timestamp 1732044439
transform 1 0 1680 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm55
timestamp 1732044439
transform 1 0 1960 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm56
timestamp 1732044439
transform 1 0 2240 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm57
timestamp 1732044439
transform 1 0 2520 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm58
timestamp 1732044439
transform 1 0 2800 0 1 -6600
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm59
timestamp 1732044439
transform 1 0 280 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm60
timestamp 1732044439
transform 1 0 560 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm61
timestamp 1732044439
transform 1 0 840 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm62
timestamp 1732044439
transform 1 0 1120 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm63
timestamp 1732044439
transform 1 0 1400 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm64
timestamp 1732044439
transform 1 0 1680 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm65
timestamp 1732044439
transform 1 0 1960 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm66
timestamp 1732044439
transform 1 0 2240 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm67
timestamp 1732044439
transform 1 0 2520 0 1 -7360
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm68
timestamp 1732044439
transform 1 0 2800 0 1 -7360
box -73 -257 73 257
<< end >>
