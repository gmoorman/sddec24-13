magic
tech sky130B
magscale 1 2
timestamp 1734220434
<< metal1 >>
rect 340 2980 540 3180
rect 920 2980 1120 3180
rect 440 80 500 2980
rect 620 2800 820 2820
rect 620 2760 640 2800
rect 630 2740 640 2760
rect 820 2740 830 2760
rect 960 720 1040 2980
rect 980 80 1040 720
rect 1220 2620 1420 2880
rect 1220 2540 1260 2620
rect 1380 2540 1420 2620
rect 1220 580 1420 2540
rect 1320 220 1420 580
rect 440 -20 520 80
rect 940 -20 1040 80
rect 540 -2000 640 -1940
rect 800 -2000 940 -1940
<< via1 >>
rect 640 2740 820 2800
rect 1260 2540 1380 2620
rect 640 -2000 800 -1940
<< metal2 >>
rect 640 2800 820 2810
rect 1220 2800 1420 2880
rect 820 2740 1420 2800
rect 640 2730 820 2740
rect 1220 2680 1420 2740
rect 1260 2620 1380 2630
rect 1260 2530 1380 2540
rect 2197 57 2404 260
rect 2199 -1078 2402 57
rect 1319 -1281 2402 -1078
rect 640 -1940 800 -1930
rect 1319 -1940 1522 -1281
rect 800 -2000 1522 -1940
rect 640 -2010 800 -2000
use inverter  x1
timestamp 1734219447
transform 1 0 1680 0 1 -820
box -360 100 720 2080
use sky130_fd_pr__nfet_g5v0d10v5_PXKL9Z  XM1
timestamp 1734219447
transform 1 0 728 0 1 1718
box -428 -1258 428 1258
use sky130_fd_pr__pfet_g5v0d10v5_V6BEPM  XM2
timestamp 1734220272
transform 1 0 738 0 1 -903
box -458 -1297 458 1297
<< labels >>
flabel metal1 340 2980 540 3180 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 920 2980 1120 3180 0 FreeSans 256 0 0 0 Vout
port 0 nsew
flabel metal2 1220 2680 1420 2880 0 FreeSans 256 0 0 0 En
port 2 nsew
<< end >>
