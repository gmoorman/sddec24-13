magic
tech sky130B
magscale 1 2
timestamp 1733700048
<< nwell >>
rect -296 -3155 296 3155
<< pmoslvt >>
rect -100 1136 100 2936
rect -100 -900 100 900
rect -100 -2936 100 -1136
<< pdiff >>
rect -158 2924 -100 2936
rect -158 1148 -146 2924
rect -112 1148 -100 2924
rect -158 1136 -100 1148
rect 100 2924 158 2936
rect 100 1148 112 2924
rect 146 1148 158 2924
rect 100 1136 158 1148
rect -158 888 -100 900
rect -158 -888 -146 888
rect -112 -888 -100 888
rect -158 -900 -100 -888
rect 100 888 158 900
rect 100 -888 112 888
rect 146 -888 158 888
rect 100 -900 158 -888
rect -158 -1148 -100 -1136
rect -158 -2924 -146 -1148
rect -112 -2924 -100 -1148
rect -158 -2936 -100 -2924
rect 100 -1148 158 -1136
rect 100 -2924 112 -1148
rect 146 -2924 158 -1148
rect 100 -2936 158 -2924
<< pdiffc >>
rect -146 1148 -112 2924
rect 112 1148 146 2924
rect -146 -888 -112 888
rect 112 -888 146 888
rect -146 -2924 -112 -1148
rect 112 -2924 146 -1148
<< nsubdiff >>
rect -260 3085 -164 3119
rect 164 3085 260 3119
rect -260 3023 -226 3085
rect 226 3023 260 3085
rect -260 -3085 -226 -3023
rect 226 -3085 260 -3023
rect -260 -3119 -164 -3085
rect 164 -3119 260 -3085
<< nsubdiffcont >>
rect -164 3085 164 3119
rect -260 -3023 -226 3023
rect 226 -3023 260 3023
rect -164 -3119 164 -3085
<< poly >>
rect -100 3017 100 3033
rect -100 2983 -84 3017
rect 84 2983 100 3017
rect -100 2936 100 2983
rect -100 1089 100 1136
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 1039 100 1055
rect -100 981 100 997
rect -100 947 -84 981
rect 84 947 100 981
rect -100 900 100 947
rect -100 -947 100 -900
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -997 100 -981
rect -100 -1055 100 -1039
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -100 -1136 100 -1089
rect -100 -2983 100 -2936
rect -100 -3017 -84 -2983
rect 84 -3017 100 -2983
rect -100 -3033 100 -3017
<< polycont >>
rect -84 2983 84 3017
rect -84 1055 84 1089
rect -84 947 84 981
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -84 -3017 84 -2983
<< locali >>
rect -260 3085 -164 3119
rect 164 3085 260 3119
rect -260 3023 -226 3085
rect 226 3023 260 3085
rect -100 2983 -84 3017
rect 84 2983 100 3017
rect -146 2924 -112 2940
rect -146 1132 -112 1148
rect 112 2924 146 2940
rect 112 1132 146 1148
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 947 -84 981
rect 84 947 100 981
rect -146 888 -112 904
rect -146 -904 -112 -888
rect 112 888 146 904
rect 112 -904 146 -888
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -146 -1148 -112 -1132
rect -146 -2940 -112 -2924
rect 112 -1148 146 -1132
rect 112 -2940 146 -2924
rect -100 -3017 -84 -2983
rect 84 -3017 100 -2983
rect -260 -3085 -226 -3023
rect 226 -3085 260 -3023
rect -260 -3119 -164 -3085
rect 164 -3119 260 -3085
<< viali >>
rect -84 2983 84 3017
rect -146 1148 -112 2924
rect 112 1148 146 2924
rect -84 1055 84 1089
rect -84 947 84 981
rect -146 -888 -112 888
rect 112 -888 146 888
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -146 -2924 -112 -1148
rect 112 -2924 146 -1148
rect -84 -3017 84 -2983
<< metal1 >>
rect -96 3017 96 3023
rect -96 2983 -84 3017
rect 84 2983 96 3017
rect -96 2977 96 2983
rect -152 2924 -106 2936
rect -152 1148 -146 2924
rect -112 1148 -106 2924
rect -152 1136 -106 1148
rect 106 2924 152 2936
rect 106 1148 112 2924
rect 146 1148 152 2924
rect 106 1136 152 1148
rect -96 1089 96 1095
rect -96 1055 -84 1089
rect 84 1055 96 1089
rect -96 1049 96 1055
rect -96 981 96 987
rect -96 947 -84 981
rect 84 947 96 981
rect -96 941 96 947
rect -152 888 -106 900
rect -152 -888 -146 888
rect -112 -888 -106 888
rect -152 -900 -106 -888
rect 106 888 152 900
rect 106 -888 112 888
rect 146 -888 152 888
rect 106 -900 152 -888
rect -96 -947 96 -941
rect -96 -981 -84 -947
rect 84 -981 96 -947
rect -96 -987 96 -981
rect -96 -1055 96 -1049
rect -96 -1089 -84 -1055
rect 84 -1089 96 -1055
rect -96 -1095 96 -1089
rect -152 -1148 -106 -1136
rect -152 -2924 -146 -1148
rect -112 -2924 -106 -1148
rect -152 -2936 -106 -2924
rect 106 -1148 152 -1136
rect 106 -2924 112 -1148
rect 146 -2924 152 -1148
rect 106 -2936 152 -2924
rect -96 -2983 96 -2977
rect -96 -3017 -84 -2983
rect 84 -3017 96 -2983
rect -96 -3023 96 -3017
<< properties >>
string FIXED_BBOX -243 -3102 243 3102
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 9.0 l 1.0 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
