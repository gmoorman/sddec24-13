magic
tech sky130B
magscale 1 2
timestamp 1733215642
<< nwell >>
rect -331 -121 1363 1163
<< nsubdiff >>
rect -295 1093 -235 1127
rect 1267 1093 1327 1127
rect -295 1067 -261 1093
rect -295 -51 -261 -25
rect 1293 1067 1327 1093
rect 1293 -51 1327 -25
rect -295 -85 -235 -51
rect 1267 -85 1327 -51
<< nsubdiffcont >>
rect -235 1093 1267 1127
rect -295 -25 -261 1067
rect 1293 -25 1327 1067
rect -235 -85 1267 -51
<< locali >>
rect -295 1093 -235 1127
rect 1267 1093 1327 1127
rect -295 1067 -261 1093
rect 1293 1067 1327 1093
rect -295 -51 -261 -25
rect 1293 -51 1327 -25
rect -295 -85 -235 -51
rect 1267 -85 1327 -51
<< viali >>
rect 1290 702 1293 796
rect 1293 702 1327 796
rect 1327 702 1328 796
<< metal1 >>
rect 556 1014 652 1030
rect 556 966 866 1014
rect 556 942 652 966
rect 1284 796 1334 808
rect 1284 770 1290 796
rect 1246 768 1290 770
rect 38 592 98 748
rect 1162 732 1290 768
rect 268 592 314 704
rect 1162 690 1206 732
rect 1246 730 1290 732
rect 1284 702 1290 730
rect 1328 702 1334 796
rect 1284 690 1334 702
rect 890 628 1016 630
rect 776 592 1016 628
rect 776 590 902 592
rect 784 444 910 482
rect 310 378 348 386
rect 342 364 490 366
rect 540 364 664 366
rect 24 360 110 362
rect 342 360 664 364
rect 24 330 664 360
rect 24 328 110 330
rect 342 328 664 330
rect 342 326 490 328
rect 632 160 664 328
rect 798 292 894 302
rect 976 292 1016 592
rect 798 254 1016 292
rect 798 214 894 254
rect 44 108 90 110
rect 608 108 704 160
rect 1164 108 1206 690
rect 44 68 1210 108
rect 44 32 90 68
rect 310 64 1210 68
use sky130_fd_pr__pfet_01v8_MJB5SZ  sky130_fd_pr__pfet_01v8_MJB5SZ_0
timestamp 1733210498
transform 1 0 287 0 1 350
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJB5SZ  sky130_fd_pr__pfet_01v8_MJB5SZ_1
timestamp 1733210498
transform 1 0 69 0 1 348
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJB5SZ  sky130_fd_pr__pfet_01v8_MJB5SZ_2
timestamp 1733210498
transform 1 0 843 0 1 724
box -109 -300 109 300
<< labels >>
rlabel metal1 798 214 894 302 1 out
port 3 n
rlabel metal1 556 942 652 1030 1 VDD
port 1 n
rlabel metal1 608 72 704 160 1 VSS
port 4 n
<< end >>
