magic
tech sky130B
timestamp 1734219447
<< pwell >>
rect -214 -629 214 629
<< mvnmos >>
rect -100 -500 100 500
<< mvndiff >>
rect -129 494 -100 500
rect -129 -494 -123 494
rect -106 -494 -100 494
rect -129 -500 -100 -494
rect 100 494 129 500
rect 100 -494 106 494
rect 123 -494 129 494
rect 100 -500 129 -494
<< mvndiffc >>
rect -123 -494 -106 494
rect 106 -494 123 494
<< mvpsubdiff >>
rect -196 605 196 611
rect -196 588 -142 605
rect 142 588 196 605
rect -196 582 196 588
rect -196 557 -167 582
rect -196 -557 -190 557
rect -173 -557 -167 557
rect 167 557 196 582
rect -196 -582 -167 -557
rect 167 -557 173 557
rect 190 -557 196 557
rect 167 -582 196 -557
rect -196 -588 196 -582
rect -196 -605 -142 -588
rect 142 -605 196 -588
rect -196 -611 196 -605
<< mvpsubdiffcont >>
rect -142 588 142 605
rect -190 -557 -173 557
rect 173 -557 190 557
rect -142 -605 142 -588
<< poly >>
rect -100 536 100 544
rect -100 519 -92 536
rect 92 519 100 536
rect -100 500 100 519
rect -100 -519 100 -500
rect -100 -536 -92 -519
rect 92 -536 100 -519
rect -100 -544 100 -536
<< polycont >>
rect -92 519 92 536
rect -92 -536 92 -519
<< locali >>
rect -190 588 -142 605
rect 142 588 190 605
rect -190 557 -173 588
rect 173 557 190 588
rect -100 519 -92 536
rect 92 519 100 536
rect -123 494 -106 502
rect -123 -502 -106 -494
rect 106 494 123 502
rect 106 -502 123 -494
rect -100 -536 -92 -519
rect 92 -536 100 -519
rect -190 -588 -173 -557
rect 173 -588 190 -557
rect -190 -605 -142 -588
rect 142 -605 190 -588
<< viali >>
rect -92 519 92 536
rect -123 -494 -106 494
rect 106 -494 123 494
rect -92 -536 92 -519
<< metal1 >>
rect -98 536 98 539
rect -98 519 -92 536
rect 92 519 98 536
rect -98 516 98 519
rect -126 494 -103 500
rect -126 -494 -123 494
rect -106 -494 -103 494
rect -126 -500 -103 -494
rect 103 494 126 500
rect 103 -494 106 494
rect 123 -494 126 494
rect 103 -500 126 -494
rect -98 -519 98 -516
rect -98 -536 -92 -519
rect 92 -536 98 -519
rect -98 -539 98 -536
<< properties >>
string FIXED_BBOX -181 -596 181 596
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
