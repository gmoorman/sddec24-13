magic
tech sky130B
magscale 1 2
timestamp 1729978887
<< nwell >>
rect -38 262 590 582
<< pwell >>
rect 0 19 552 159
rect 29 -17 63 19
<< nmos >>
rect 149 47 179 131
rect 373 47 403 131
<< pmos >>
rect 149 413 179 497
rect 373 413 403 497
<< ndiff >>
rect 27 106 149 131
rect 27 72 35 106
rect 69 72 149 106
rect 27 47 149 72
rect 179 47 373 131
rect 403 106 525 131
rect 403 72 483 106
rect 517 72 525 106
rect 403 47 525 72
<< pdiff >>
rect 27 472 149 497
rect 27 438 35 472
rect 69 438 149 472
rect 27 413 149 438
rect 179 472 373 497
rect 179 438 259 472
rect 293 438 373 472
rect 179 413 373 438
rect 403 472 525 497
rect 403 438 483 472
rect 517 438 525 472
rect 403 413 525 438
<< ndiffc >>
rect 35 72 69 106
rect 483 72 517 106
<< pdiffc >>
rect 35 438 69 472
rect 259 438 293 472
rect 483 438 517 472
<< poly >>
rect 149 497 179 523
rect 373 497 403 523
rect 149 312 179 413
rect 84 297 179 312
rect 84 263 121 297
rect 155 263 179 297
rect 373 272 403 413
rect 84 232 179 263
rect 149 131 179 232
rect 308 253 403 272
rect 308 219 327 253
rect 361 219 403 253
rect 308 192 403 219
rect 373 131 403 192
rect 149 21 179 47
rect 373 21 403 47
<< polycont >>
rect 121 263 155 297
rect 327 219 361 253
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 35 472 69 527
rect 35 421 69 438
rect 259 472 293 489
rect 259 349 293 438
rect 483 472 517 527
rect 483 421 517 438
rect 259 332 517 349
rect 96 297 176 330
rect 259 315 523 332
rect 96 263 121 297
rect 155 263 176 297
rect 96 260 176 263
rect 294 253 380 270
rect 294 219 327 253
rect 361 219 380 253
rect 294 208 380 219
rect 460 212 523 315
rect 35 106 69 123
rect 35 17 69 72
rect 483 106 517 212
rect 483 55 517 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel nwell 29 527 63 561 0 FreeSans 240 0 0 0 VPB
port 1 nsew power bidirectional
flabel metal1 29 527 63 561 0 FreeSans 240 0 0 0 VPWR
port 2 nsew
flabel pwell 29 -17 63 17 0 FreeSans 240 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 29 -17 63 17 0 FreeSans 240 0 0 0 VGND
port 4 nsew
flabel locali 121 289 155 323 0 FreeSans 240 0 0 0 A
port 5 nsew signal input
flabel locali 305 221 339 255 0 FreeSans 240 0 0 0 B
port 6 nsew signal output
flabel locali 489 289 523 323 0 FreeSans 240 0 0 0 X
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 552 544
<< end >>
