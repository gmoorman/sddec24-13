magic
tech sky130B
magscale 1 2
timestamp 1733717322
<< xpolycontact >>
rect -573 7526 573 7958
rect -573 6994 573 7426
rect -573 6458 573 6890
rect -573 5926 573 6358
rect -573 5390 573 5822
rect -573 4858 573 5290
rect -573 4322 573 4754
rect -573 3790 573 4222
rect -573 3254 573 3686
rect -573 2722 573 3154
rect -573 2186 573 2618
rect -573 1654 573 2086
rect -573 1118 573 1550
rect -573 586 573 1018
rect -573 50 573 482
rect -573 -482 573 -50
rect -573 -1018 573 -586
rect -573 -1550 573 -1118
rect -573 -2086 573 -1654
rect -573 -2618 573 -2186
rect -573 -3154 573 -2722
rect -573 -3686 573 -3254
rect -573 -4222 573 -3790
rect -573 -4754 573 -4322
rect -573 -5290 573 -4858
rect -573 -5822 573 -5390
rect -573 -6358 573 -5926
rect -573 -6890 573 -6458
rect -573 -7426 573 -6994
rect -573 -7958 573 -7526
<< ppolyres >>
rect -573 7426 573 7526
rect -573 6358 573 6458
rect -573 5290 573 5390
rect -573 4222 573 4322
rect -573 3154 573 3254
rect -573 2086 573 2186
rect -573 1018 573 1118
rect -573 -50 573 50
rect -573 -1118 573 -1018
rect -573 -2186 573 -2086
rect -573 -3254 573 -3154
rect -573 -4322 573 -4222
rect -573 -5390 573 -5290
rect -573 -6458 573 -6358
rect -573 -7526 573 -7426
<< viali >>
rect -557 7543 557 7940
rect -557 7012 557 7409
rect -557 6475 557 6872
rect -557 5944 557 6341
rect -557 5407 557 5804
rect -557 4876 557 5273
rect -557 4339 557 4736
rect -557 3808 557 4205
rect -557 3271 557 3668
rect -557 2740 557 3137
rect -557 2203 557 2600
rect -557 1672 557 2069
rect -557 1135 557 1532
rect -557 604 557 1001
rect -557 67 557 464
rect -557 -464 557 -67
rect -557 -1001 557 -604
rect -557 -1532 557 -1135
rect -557 -2069 557 -1672
rect -557 -2600 557 -2203
rect -557 -3137 557 -2740
rect -557 -3668 557 -3271
rect -557 -4205 557 -3808
rect -557 -4736 557 -4339
rect -557 -5273 557 -4876
rect -557 -5804 557 -5407
rect -557 -6341 557 -5944
rect -557 -6872 557 -6475
rect -557 -7409 557 -7012
rect -557 -7940 557 -7543
<< metal1 >>
rect -569 7940 569 7946
rect -569 7543 -557 7940
rect 557 7543 569 7940
rect -569 7537 569 7543
rect -569 7409 569 7415
rect -569 7012 -557 7409
rect 557 7012 569 7409
rect -569 7006 569 7012
rect -569 6872 569 6878
rect -569 6475 -557 6872
rect 557 6475 569 6872
rect -569 6469 569 6475
rect -569 6341 569 6347
rect -569 5944 -557 6341
rect 557 5944 569 6341
rect -569 5938 569 5944
rect -569 5804 569 5810
rect -569 5407 -557 5804
rect 557 5407 569 5804
rect -569 5401 569 5407
rect -569 5273 569 5279
rect -569 4876 -557 5273
rect 557 4876 569 5273
rect -569 4870 569 4876
rect -569 4736 569 4742
rect -569 4339 -557 4736
rect 557 4339 569 4736
rect -569 4333 569 4339
rect -569 4205 569 4211
rect -569 3808 -557 4205
rect 557 3808 569 4205
rect -569 3802 569 3808
rect -569 3668 569 3674
rect -569 3271 -557 3668
rect 557 3271 569 3668
rect -569 3265 569 3271
rect -569 3137 569 3143
rect -569 2740 -557 3137
rect 557 2740 569 3137
rect -569 2734 569 2740
rect -569 2600 569 2606
rect -569 2203 -557 2600
rect 557 2203 569 2600
rect -569 2197 569 2203
rect -569 2069 569 2075
rect -569 1672 -557 2069
rect 557 1672 569 2069
rect -569 1666 569 1672
rect -569 1532 569 1538
rect -569 1135 -557 1532
rect 557 1135 569 1532
rect -569 1129 569 1135
rect -569 1001 569 1007
rect -569 604 -557 1001
rect 557 604 569 1001
rect -569 598 569 604
rect -569 464 569 470
rect -569 67 -557 464
rect 557 67 569 464
rect -569 61 569 67
rect -569 -67 569 -61
rect -569 -464 -557 -67
rect 557 -464 569 -67
rect -569 -470 569 -464
rect -569 -604 569 -598
rect -569 -1001 -557 -604
rect 557 -1001 569 -604
rect -569 -1007 569 -1001
rect -569 -1135 569 -1129
rect -569 -1532 -557 -1135
rect 557 -1532 569 -1135
rect -569 -1538 569 -1532
rect -569 -1672 569 -1666
rect -569 -2069 -557 -1672
rect 557 -2069 569 -1672
rect -569 -2075 569 -2069
rect -569 -2203 569 -2197
rect -569 -2600 -557 -2203
rect 557 -2600 569 -2203
rect -569 -2606 569 -2600
rect -569 -2740 569 -2734
rect -569 -3137 -557 -2740
rect 557 -3137 569 -2740
rect -569 -3143 569 -3137
rect -569 -3271 569 -3265
rect -569 -3668 -557 -3271
rect 557 -3668 569 -3271
rect -569 -3674 569 -3668
rect -569 -3808 569 -3802
rect -569 -4205 -557 -3808
rect 557 -4205 569 -3808
rect -569 -4211 569 -4205
rect -569 -4339 569 -4333
rect -569 -4736 -557 -4339
rect 557 -4736 569 -4339
rect -569 -4742 569 -4736
rect -569 -4876 569 -4870
rect -569 -5273 -557 -4876
rect 557 -5273 569 -4876
rect -569 -5279 569 -5273
rect -569 -5407 569 -5401
rect -569 -5804 -557 -5407
rect 557 -5804 569 -5407
rect -569 -5810 569 -5804
rect -569 -5944 569 -5938
rect -569 -6341 -557 -5944
rect 557 -6341 569 -5944
rect -569 -6347 569 -6341
rect -569 -6475 569 -6469
rect -569 -6872 -557 -6475
rect 557 -6872 569 -6475
rect -569 -6878 569 -6872
rect -569 -7012 569 -7006
rect -569 -7409 -557 -7012
rect 557 -7409 569 -7012
rect -569 -7415 569 -7409
rect -569 -7543 569 -7537
rect -569 -7940 -557 -7543
rect 557 -7940 569 -7543
rect -569 -7946 569 -7940
<< properties >>
string gencell sky130_fd_pr__res_high_po_5p73
string library sky130
string parameters w 5.730 l 0.5 m 15 nx 1 wmin 5.730 lmin 0.50 rho 319.8 val 1.099k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 1 full_metal 0 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
