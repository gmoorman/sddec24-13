** sch_path: /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/xschem/userLib/4bitADC.sch
**.subckt 4bitADC
R1 net1 Vrefa sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R2 net2 net1 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
x1 VDD net3 net22 Clk Vin net1 GND Comparator
R3 net4 net2 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R4 net5 net4 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R5 net6 net5 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R6 net7 net6 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R7 net8 net7 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R8 net9 net8 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R9 net10 net9 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R10 GND net10 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
V1 VDD GND 5
V2 Clk GND pulse(0 5 1ns 1ns 1ns 500ns 1us)
V3 Vrefa GND 5
V4 Vin GND sin(2.5 2.5 100k)
x3 VDD net11 net23 Clk Vin net4 GND Comparator
x5 VDD net12 net24 Clk Vin net6 GND Comparator
x7 VDD net13 net25 Clk Vin net8 GND Comparator
x9 VDD net14 net26 Clk Vin net10 GND Comparator
XM5 b3 net21 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 b3 net15 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 b2 net20 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 b2 net16 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 b1 net20 GND net18 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 b1 net16 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 b0 net21 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 b0 net20 GND net19 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R11 b3 net17 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R12 b2 net17 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R13 b1 net17 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
R14 b0 net17 sky130_fd_pr__res_generic_l1 W=1 L=5 m=1
x8 net21 net3 net11 VDD GND VDD GND AND2I
x2 net15 net11 net12 VDD GND VDD GND AND2I
x4 net20 net12 net13 VDD GND VDD GND AND2I
x6 net16 net13 net14 VDD GND VDD GND AND2I
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice



.tran 100n 10u
.save all


**** end user architecture code
**.ends

* expanding   symbol:  dependencies/pdks/sky130B/libs.tech/xschem/userLib/Comparator.sym # of pins=7
** sym_path: /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/xschem/userLib/Comparator.sym
** sch_path: /home/gmoorman/caravel_user_project/dependencies/pdks/sky130B/libs.tech/xschem/userLib/Comparator.sch
.subckt Comparator VDD V1 V2 CLK VIN VREF VSS
*.iopin VDD
*.iopin VSS
*.ipin VIN
*.ipin VREF
*.opin V2
*.opin V1
*.ipin CLK
XM7 V2 V1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.72 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 V2 CLK VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.72 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 V1 CLK VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.72 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 V1 V2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.72 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 V2 CLK net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.72 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 V1 CLK net4 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.72 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net4 V2 net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.72 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 V1 net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.72 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.72 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 VREF VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.72 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
