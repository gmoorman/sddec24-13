magic
tech sky130B
magscale 1 2
timestamp 1735082180
<< nwell >>
rect -1116 9486 37204 9588
rect -1526 9356 -728 9438
<< pwell >>
rect 13156 50 13186 6572
rect 26314 50 26344 6572
rect -4388 -186 -4358 -76
rect -1486 -186 -1446 -44
rect -454 -52 37866 50
rect -2 -186 28 -76
rect 2900 -186 2940 -52
rect 7286 -186 7326 -52
rect 11672 -186 11712 -52
rect 13156 -186 13186 -52
rect 16058 -186 16098 -52
rect 20444 -186 20484 -52
rect 24830 -186 24870 -52
rect 26314 -186 26344 -52
rect 29216 -186 29256 -52
rect 33602 -186 33642 -52
rect 37988 -186 38028 -44
rect 39472 -186 39502 6572
rect 42374 -186 42414 -44
rect 46760 -186 46800 -44
rect 51146 -186 51186 -46
rect 52630 -186 52660 6570
rect 61550 2214 61620 2268
rect 55532 -186 55572 -46
rect 59942 -186 59982 -46
rect 64300 -186 64340 -48
<< metal1 >>
rect -1116 9486 65598 9588
<< metal2 >>
rect -1264 9854 -1254 9926
rect -1182 9854 -1172 9926
rect 3122 9854 3132 9926
rect 3204 9854 3214 9926
rect 7508 9856 7518 9928
rect 7590 9856 7600 9928
rect 11894 9856 11904 9928
rect 11976 9856 11986 9928
rect 16280 9852 16290 9924
rect 16362 9852 16372 9924
rect 20668 9868 20678 9940
rect 20750 9868 20760 9940
rect 25052 9856 25062 9928
rect 25134 9856 25144 9928
rect 35926 9926 38290 9928
rect 29438 9852 29448 9924
rect 29520 9852 29530 9924
rect 34222 9906 34232 9922
rect 33888 9850 34232 9906
rect 34304 9850 34314 9922
rect 35834 9854 35844 9926
rect 35916 9856 38290 9926
rect 35916 9854 35926 9856
rect 40286 9848 40296 9920
rect 40368 9848 42692 9920
rect 46980 9854 46990 9926
rect 47062 9854 47072 9926
rect 51368 9856 51378 9928
rect 51450 9856 51460 9928
rect 55754 9850 55764 9922
rect 55836 9850 55846 9922
rect 60142 9850 60152 9922
rect 60224 9850 60234 9922
rect 64526 9850 64536 9922
rect 64608 9850 64618 9922
rect -1032 6660 -960 6670
rect -1032 6578 -960 6588
rect 3354 6662 3426 6672
rect 3354 6580 3426 6590
rect 7744 6662 7816 6672
rect 7744 6580 7816 6590
rect 12130 6662 12202 6672
rect 12130 6580 12202 6590
rect 16514 6658 16586 6668
rect 16514 6576 16586 6586
rect 20900 6662 20972 6672
rect 20900 6580 20972 6590
rect 25284 6660 25356 6670
rect 25284 6578 25356 6588
rect 29672 6662 29744 6672
rect 29672 6580 29744 6590
rect 34058 6660 34130 6670
rect 34058 6578 34130 6588
rect 38444 6662 38516 6672
rect 38444 6580 38516 6590
rect 42830 6660 42902 6670
rect 42830 6578 42902 6588
rect 47216 6658 47288 6668
rect 47216 6576 47288 6586
rect 51602 6660 51674 6670
rect 51602 6578 51674 6588
rect 55988 6662 56060 6672
rect 55988 6580 56060 6590
rect 60372 6658 60444 6668
rect 60372 6576 60444 6586
rect 64760 6658 64832 6668
rect 64760 6576 64832 6586
<< via2 >>
rect -1254 9854 -1182 9926
rect 3132 9854 3204 9926
rect 7518 9856 7590 9928
rect 11904 9856 11976 9928
rect 16290 9852 16362 9924
rect 20678 9868 20750 9940
rect 25062 9856 25134 9928
rect 29448 9852 29520 9924
rect 34232 9850 34304 9922
rect 35844 9854 35916 9926
rect 40296 9848 40368 9920
rect 46990 9854 47062 9926
rect 51378 9856 51450 9928
rect 55764 9850 55836 9922
rect 60152 9850 60224 9922
rect 64536 9850 64608 9922
rect -1032 6588 -960 6660
rect 3354 6590 3426 6662
rect 7744 6590 7816 6662
rect 12130 6590 12202 6662
rect 16514 6586 16586 6658
rect 20900 6590 20972 6662
rect 25284 6588 25356 6660
rect 29672 6590 29744 6662
rect 34058 6588 34130 6660
rect 38444 6590 38516 6662
rect 42830 6588 42902 6660
rect 47216 6586 47288 6658
rect 51602 6588 51674 6660
rect 55988 6590 56060 6662
rect 60372 6586 60444 6658
rect 64760 6586 64832 6658
<< metal3 >>
rect 32996 11810 33028 11928
rect 32996 10904 33058 11810
rect 33784 11594 33820 11714
rect -1254 10844 33058 10904
rect -1254 9936 -1180 10844
rect 33210 10784 33272 11108
rect 3118 10724 33272 10784
rect 3132 9936 3204 10724
rect 33482 10664 33544 11110
rect 7504 10604 33544 10664
rect 7518 9938 7590 10604
rect 33754 10542 33820 11594
rect 11892 10482 33820 10542
rect 11904 9938 11976 10482
rect 34026 10422 34092 11108
rect 16276 10362 34094 10422
rect -1259 9926 -1177 9936
rect -1259 9854 -1254 9926
rect -1182 9854 -1177 9926
rect -1259 9844 -1177 9854
rect 3127 9926 3209 9936
rect 3127 9854 3132 9926
rect 3204 9854 3209 9926
rect 3127 9844 3209 9854
rect 7513 9928 7595 9938
rect 7513 9856 7518 9928
rect 7590 9856 7595 9928
rect 7513 9846 7595 9856
rect 11899 9928 11981 9938
rect 16290 9934 16362 10362
rect 20678 10300 34112 10302
rect 34294 10300 34360 11116
rect 20678 10238 34360 10300
rect 20678 9950 20750 10238
rect 34570 10178 34636 11116
rect 25042 10118 34636 10178
rect 20673 9940 20755 9950
rect 11899 9856 11904 9928
rect 11976 9856 11981 9928
rect 11899 9846 11981 9856
rect 16285 9924 16367 9934
rect 16285 9852 16290 9924
rect 16362 9852 16367 9924
rect 20673 9868 20678 9940
rect 20750 9868 20755 9940
rect 25062 9938 25142 10118
rect 34840 10058 34906 11116
rect 29434 9998 34906 10058
rect 35110 10874 35176 11110
rect 35430 10878 35496 11116
rect 35700 10878 35766 11118
rect 35980 10880 36046 11110
rect 36252 10882 36318 11110
rect 36524 10882 36590 11110
rect 29434 9994 34640 9998
rect 20673 9858 20755 9868
rect 25057 9928 25142 9938
rect 16285 9842 16367 9852
rect 25057 9856 25062 9928
rect 25134 9858 25142 9928
rect 29442 9924 29526 9994
rect 25134 9856 25139 9858
rect 25057 9846 25139 9856
rect 29442 9854 29448 9924
rect 29443 9852 29448 9854
rect 29520 9854 29526 9924
rect 34227 9922 34309 9932
rect 29520 9852 29525 9854
rect 29443 9842 29525 9852
rect 34227 9850 34232 9922
rect 34304 9850 34309 9922
rect 34227 9840 34309 9850
rect 34230 9780 34308 9840
rect 34230 9778 34958 9780
rect 35110 9778 35178 10874
rect 35430 9784 35506 10878
rect 35700 10056 35776 10878
rect 35980 10176 36050 10880
rect 36252 10302 36322 10882
rect 36524 10424 36594 10882
rect 36796 10546 36866 11062
rect 37072 10670 37142 11068
rect 37072 10668 37898 10670
rect 37072 10608 64640 10668
rect 36796 10544 37622 10546
rect 36796 10484 60236 10544
rect 36524 10422 37350 10424
rect 36524 10362 55836 10422
rect 36252 10296 37058 10302
rect 36252 10236 51460 10296
rect 51062 10234 51460 10236
rect 35980 10116 47074 10176
rect 35700 9996 40368 10056
rect 35839 9926 35921 9936
rect 40296 9930 40368 9996
rect 46990 9936 47060 10116
rect 51376 9938 51460 10234
rect 35839 9854 35844 9926
rect 35916 9854 35921 9926
rect 35839 9844 35921 9854
rect 40291 9920 40373 9930
rect 40291 9848 40296 9920
rect 40368 9848 40373 9920
rect 35842 9784 35916 9844
rect 40291 9838 40373 9848
rect 46985 9926 47067 9936
rect 46985 9854 46990 9926
rect 47062 9854 47067 9926
rect 46985 9844 47067 9854
rect 51373 9928 51460 9938
rect 55764 9932 55836 10362
rect 60152 9932 60236 10484
rect 64536 9932 64612 10608
rect 51373 9856 51378 9928
rect 51450 9856 51460 9928
rect 55759 9922 55841 9932
rect 51373 9846 51455 9856
rect 55759 9850 55764 9922
rect 55836 9850 55841 9922
rect 55759 9840 55841 9850
rect 60147 9922 60236 9932
rect 60147 9850 60152 9922
rect 60224 9850 60236 9922
rect 64531 9922 64613 9932
rect 64531 9850 64536 9922
rect 64608 9850 64613 9922
rect 60147 9840 60229 9850
rect 64531 9840 64613 9850
rect 34230 9718 35176 9778
rect 35430 9720 35920 9784
rect -1042 6660 -950 6665
rect 3344 6662 3436 6667
rect -1042 6658 -1032 6660
rect -4742 6588 -1032 6658
rect -960 6658 -898 6660
rect 3344 6658 3354 6662
rect -960 6590 3354 6658
rect 3426 6658 3436 6662
rect 7734 6662 7826 6667
rect 7734 6658 7744 6662
rect 3426 6590 7744 6658
rect 7816 6658 7826 6662
rect 12120 6662 12212 6667
rect 12120 6658 12130 6662
rect 7816 6590 12130 6658
rect 12202 6658 12212 6662
rect 16504 6658 16596 6663
rect 20890 6662 20982 6667
rect 20890 6658 20900 6662
rect 12202 6590 16514 6658
rect -960 6588 16514 6590
rect -4742 6586 16514 6588
rect 16586 6590 20900 6658
rect 20972 6658 20982 6662
rect 25274 6660 25366 6665
rect 25274 6658 25284 6660
rect 20972 6590 25284 6658
rect 16586 6588 25284 6590
rect 25356 6658 25366 6660
rect 29662 6662 29754 6667
rect 29662 6658 29672 6662
rect 25356 6590 29672 6658
rect 29744 6658 29754 6662
rect 34048 6660 34140 6665
rect 34048 6658 34058 6660
rect 29744 6590 34058 6658
rect 25356 6588 34058 6590
rect 34130 6658 34140 6660
rect 38434 6662 38526 6667
rect 38434 6658 38444 6662
rect 34130 6590 38444 6658
rect 38516 6658 38526 6662
rect 42820 6660 42912 6665
rect 42820 6658 42830 6660
rect 38516 6590 42830 6658
rect 34130 6588 42830 6590
rect 42902 6658 42912 6660
rect 47206 6658 47298 6663
rect 51592 6660 51684 6665
rect 51592 6658 51602 6660
rect 42902 6588 47216 6658
rect 16586 6586 47216 6588
rect 47288 6588 51602 6658
rect 51674 6658 51684 6660
rect 55978 6662 56070 6667
rect 55978 6658 55988 6662
rect 51674 6590 55988 6658
rect 56060 6658 56070 6662
rect 60362 6658 60454 6663
rect 64750 6658 64842 6663
rect 56060 6590 60372 6658
rect 51674 6588 60372 6590
rect 47288 6586 60372 6588
rect 60444 6586 64760 6658
rect 64832 6586 64842 6658
rect -1042 6583 -950 6586
rect 3344 6585 3436 6586
rect 7734 6585 7826 6586
rect 12120 6585 12212 6586
rect 16504 6581 16596 6586
rect 20890 6585 20982 6586
rect 25274 6583 25366 6586
rect 29662 6585 29754 6586
rect 34048 6583 34140 6586
rect 38434 6585 38526 6586
rect 42820 6583 42912 6586
rect 47206 6581 47298 6586
rect 51592 6583 51684 6586
rect 55978 6585 56070 6586
rect 60362 6581 60454 6586
rect 64750 6581 64842 6586
use combination_test_DUMMY  combination_test_DUMMY_0
timestamp 1733627311
transform 1 0 53078 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_1
timestamp 1733627311
transform 1 0 446 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_2
timestamp 1733627311
transform 1 0 39920 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_3
timestamp 1733627311
transform 1 0 48692 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_4
timestamp 1733627311
transform 1 0 44306 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_5
timestamp 1733627311
transform 1 0 17990 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_6
timestamp 1733627311
transform 1 0 13604 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_7
timestamp 1733627311
transform 1 0 9218 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_8
timestamp 1733627311
transform 1 0 4832 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_9
timestamp 1733627311
transform 1 0 22376 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_10
timestamp 1733627311
transform 1 0 26762 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_11
timestamp 1733627311
transform 1 0 31148 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_12
timestamp 1733627311
transform 1 0 35534 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_13
timestamp 1733627311
transform 1 0 57464 0 1 8470
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_14
timestamp 1733627311
transform 1 0 61850 0 1 8470
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_15
timestamp 1733627311
transform 1 0 -3940 0 1 8472
box -574 -8600 3812 1466
use Priority_Encoder_16t4  Priority_Encoder_16t4_1
timestamp 1733718626
transform 0 -1 39060 -1 0 19032
box 0 1096 8000 6928
<< end >>
