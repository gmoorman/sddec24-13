magic
tech sky130B
magscale 1 2
timestamp 1729979448
<< error_s >>
rect 298 4915 333 4949
rect 299 4896 333 4915
rect 129 4847 187 4853
rect 129 4813 141 4847
rect 129 4807 187 4813
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 4896
rect 352 4862 387 4896
rect 352 583 386 4862
rect 498 4794 556 4800
rect 498 4760 510 4794
rect 498 4754 556 4760
rect 1774 4685 1809 4719
rect 1775 4666 1809 4685
rect 1605 4617 1663 4623
rect 1605 4583 1617 4617
rect 1605 4577 1663 4583
rect 668 1643 702 1697
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 687 530 702 1643
rect 721 1609 756 1643
rect 1036 1609 1071 1643
rect 1459 1626 1493 1644
rect 721 530 755 1609
rect 1037 1590 1071 1609
rect 867 1541 925 1547
rect 867 1507 879 1541
rect 867 1501 925 1507
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1056 477 1071 1590
rect 1090 1556 1125 1590
rect 1090 477 1124 1556
rect 1236 1488 1294 1494
rect 1236 1454 1248 1488
rect 1236 1448 1294 1454
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1423 424 1493 1626
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1794 371 1809 4666
rect 1828 4632 1863 4666
rect 1828 371 1862 4632
rect 1974 4564 2032 4570
rect 1974 4530 1986 4564
rect 1974 4524 2032 4530
rect 3250 2473 3285 2507
rect 3251 2454 3285 2473
rect 3081 2405 3139 2411
rect 3081 2371 3093 2405
rect 3081 2365 3139 2371
rect 2144 1413 2178 1467
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2163 318 2178 1413
rect 2197 1379 2232 1413
rect 2512 1379 2547 1413
rect 2197 318 2231 1379
rect 2513 1360 2547 1379
rect 2343 1311 2401 1317
rect 2343 1277 2355 1311
rect 2343 1271 2401 1277
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2532 265 2547 1360
rect 2566 1326 2601 1360
rect 2566 265 2600 1326
rect 2712 1258 2770 1264
rect 2712 1224 2724 1258
rect 2712 1218 2770 1224
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect 2901 212 2916 1360
rect 2935 212 2969 1414
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3270 159 3285 2454
rect 3304 2420 3339 2454
rect 3304 159 3338 2420
rect 3450 2352 3508 2358
rect 3450 2318 3462 2352
rect 3450 2312 3508 2318
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 2454
rect 3673 106 3707 2508
rect 3673 72 3688 106
rect 3769 53 4097 87
rect 3915 0 3949 53
rect 4755 -519 4779 -495
rect 3891 -553 3915 -529
rect 4779 -543 4803 -519
rect 3915 -577 3939 -553
rect 4721 -981 4745 -957
rect 4779 -981 4803 -957
rect 4745 -1005 4779 -981
<< psubdiffcont >>
rect 3915 -519 3949 87
rect 3915 -553 4779 -519
rect 4745 -981 4779 -553
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use sky130_fd_pr__pfet_01v8_K4JMRH  XM1
timestamp 1729978744
transform 1 0 158 0 1 2766
box -211 -2219 211 2219
use sky130_fd_pr__pfet_01v8_K4JMRH  XM2
timestamp 1729978744
transform 1 0 527 0 1 2713
box -211 -2219 211 2219
use sky130_fd_pr__pfet_01v8_Y4MTK2  XM3
timestamp 1729978744
transform 1 0 896 0 1 1060
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_Y4MTK2  XM4
timestamp 1729978744
transform 1 0 1265 0 1 1007
box -211 -619 211 619
use sky130_fd_pr__nfet_01v8_NZEYJE  XM5
timestamp 1729978744
transform 1 0 1634 0 1 2545
box -211 -2210 211 2210
use sky130_fd_pr__nfet_01v8_NZEYJE  XM6
timestamp 1729978744
transform 1 0 2003 0 1 2492
box -211 -2210 211 2210
use sky130_fd_pr__nfet_01v8_N5NU4P  XM7
timestamp 1729978744
transform 1 0 2372 0 1 839
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_N5NU4P  XM8
timestamp 1729978744
transform 1 0 2741 0 1 786
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_6SJULU  XM9
timestamp 1729978744
transform 1 0 3110 0 1 1333
box -211 -1210 211 1210
use sky130_fd_pr__nfet_01v8_6SJULU  XM10
timestamp 1729978744
transform 1 0 3479 0 1 1280
box -211 -1210 211 1210
use sky130_fd_pr__nfet_01v8_33QZKN  XM11
timestamp 1729978744
transform 1 0 3933 0 1 2227
box -296 -2210 296 2210
use sky130_fd_pr__nfet_01v8_33QZKN  XM12
timestamp 1729978744
transform 1 0 6576 0 1 2316
box -296 -2210 296 2210
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vinplus
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vinminus
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLK
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Voutplus
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Voutminus
port 6 nsew
<< end >>
