magic
tech sky130B
magscale 1 2
timestamp 1733700048
<< metal4 >>
rect -1049 3439 1049 3480
rect -1049 1961 793 3439
rect 1029 1961 1049 3439
rect -1049 1920 1049 1961
rect -1049 1639 1049 1680
rect -1049 161 793 1639
rect 1029 161 1049 1639
rect -1049 120 1049 161
rect -1049 -161 1049 -120
rect -1049 -1639 793 -161
rect 1029 -1639 1049 -161
rect -1049 -1680 1049 -1639
rect -1049 -1961 1049 -1920
rect -1049 -3439 793 -1961
rect 1029 -3439 1049 -1961
rect -1049 -3480 1049 -3439
<< via4 >>
rect 793 1961 1029 3439
rect 793 161 1029 1639
rect 793 -1639 1029 -161
rect 793 -3439 1029 -1961
<< mimcap2 >>
rect -969 3360 431 3400
rect -969 2040 -929 3360
rect 391 2040 431 3360
rect -969 2000 431 2040
rect -969 1560 431 1600
rect -969 240 -929 1560
rect 391 240 431 1560
rect -969 200 431 240
rect -969 -240 431 -200
rect -969 -1560 -929 -240
rect 391 -1560 431 -240
rect -969 -1600 431 -1560
rect -969 -2040 431 -2000
rect -969 -3360 -929 -2040
rect 391 -3360 431 -2040
rect -969 -3400 431 -3360
<< mimcap2contact >>
rect -929 2040 391 3360
rect -929 240 391 1560
rect -929 -1560 391 -240
rect -929 -3360 391 -2040
<< metal5 >>
rect -429 3384 -109 3600
rect 751 3439 1071 3600
rect -953 3360 415 3384
rect -953 2040 -929 3360
rect 391 2040 415 3360
rect -953 2016 415 2040
rect -429 1584 -109 2016
rect 751 1961 793 3439
rect 1029 1961 1071 3439
rect 751 1639 1071 1961
rect -953 1560 415 1584
rect -953 240 -929 1560
rect 391 240 415 1560
rect -953 216 415 240
rect -429 -216 -109 216
rect 751 161 793 1639
rect 1029 161 1071 1639
rect 751 -161 1071 161
rect -953 -240 415 -216
rect -953 -1560 -929 -240
rect 391 -1560 415 -240
rect -953 -1584 415 -1560
rect -429 -2016 -109 -1584
rect 751 -1639 793 -161
rect 1029 -1639 1071 -161
rect 751 -1961 1071 -1639
rect -953 -2040 415 -2016
rect -953 -3360 -929 -2040
rect 391 -3360 415 -2040
rect -953 -3384 415 -3360
rect -429 -3600 -109 -3384
rect 751 -3439 793 -1961
rect 1029 -3439 1071 -1961
rect 751 -3600 1071 -3439
<< properties >>
string FIXED_BBOX -1049 1920 511 3480
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 7.0 l 7.0 val 103.32 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
