** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/4x4crossbar.sch
.subckt 4x4crossbar BL1 BL2 SL2 SL1 BL3 BL4 SL4 SL3 WL2 WL1 WL4 WL3 VSS
*.PININFO BL1:B BL2:B SL2:B SL1:B BL3:B BL4:B SL4:B SL3:B WL2:B WL1:B WL4:B WL3:B VSS:B
x1 VSS BL2 BL1 WL1 WL2 SL2 SL1 2x2crossbar
x2 VSS BL2 BL1 WL3 WL4 SL2 SL1 2x2crossbar
x3 VSS BL4 BL3 WL1 WL2 SL4 SL3 2x2crossbar
x4 VSS BL4 BL3 WL3 WL4 SL4 SL3 2x2crossbar
.ends

* expanding   symbol:  2x2crossbar.sym # of pins=7
** sym_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/2x2crossbar.sym
** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/2x2crossbar.sch
.subckt 2x2crossbar VSS BL2 BL1 WL1 WL2 SL2 SL1
*.PININFO BL2:B BL1:B VSS:B WL1:B WL2:B SL1:B SL2:B
x1 BL1 WL1 VSS SL1 1T1R
x2 BL2 WL1 VSS SL2 1T1R
x3 BL1 WL2 VSS SL1 1T1R
x4 BL2 WL2 VSS SL2 1T1R
.ends


* expanding   symbol:  1T1R.sym # of pins=4
** sym_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/1T1R.sym
** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/1T1R.sch
.subckt 1T1R BL WL VSS SL
*.PININFO SL:B VSS:B WL:B BL:B
XR1 BL net1 sky130_fd_pr_reram__reram_cell Tfilament_0=3.8e-9 area_ox=1
XM1 net1 WL SL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=1
.ends


.end
