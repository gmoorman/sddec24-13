magic
tech sky130B
magscale 1 2
timestamp 1733700048
<< nwell >>
rect -296 -2855 296 2855
<< pmoslvt >>
rect -100 1036 100 2636
rect -100 -800 100 800
rect -100 -2636 100 -1036
<< pdiff >>
rect -158 2624 -100 2636
rect -158 1048 -146 2624
rect -112 1048 -100 2624
rect -158 1036 -100 1048
rect 100 2624 158 2636
rect 100 1048 112 2624
rect 146 1048 158 2624
rect 100 1036 158 1048
rect -158 788 -100 800
rect -158 -788 -146 788
rect -112 -788 -100 788
rect -158 -800 -100 -788
rect 100 788 158 800
rect 100 -788 112 788
rect 146 -788 158 788
rect 100 -800 158 -788
rect -158 -1048 -100 -1036
rect -158 -2624 -146 -1048
rect -112 -2624 -100 -1048
rect -158 -2636 -100 -2624
rect 100 -1048 158 -1036
rect 100 -2624 112 -1048
rect 146 -2624 158 -1048
rect 100 -2636 158 -2624
<< pdiffc >>
rect -146 1048 -112 2624
rect 112 1048 146 2624
rect -146 -788 -112 788
rect 112 -788 146 788
rect -146 -2624 -112 -1048
rect 112 -2624 146 -1048
<< nsubdiff >>
rect -260 2785 -164 2819
rect 164 2785 260 2819
rect -260 2723 -226 2785
rect 226 2723 260 2785
rect -260 -2785 -226 -2723
rect 226 -2785 260 -2723
rect -260 -2819 -164 -2785
rect 164 -2819 260 -2785
<< nsubdiffcont >>
rect -164 2785 164 2819
rect -260 -2723 -226 2723
rect 226 -2723 260 2723
rect -164 -2819 164 -2785
<< poly >>
rect -100 2717 100 2733
rect -100 2683 -84 2717
rect 84 2683 100 2717
rect -100 2636 100 2683
rect -100 989 100 1036
rect -100 955 -84 989
rect 84 955 100 989
rect -100 939 100 955
rect -100 881 100 897
rect -100 847 -84 881
rect 84 847 100 881
rect -100 800 100 847
rect -100 -847 100 -800
rect -100 -881 -84 -847
rect 84 -881 100 -847
rect -100 -897 100 -881
rect -100 -955 100 -939
rect -100 -989 -84 -955
rect 84 -989 100 -955
rect -100 -1036 100 -989
rect -100 -2683 100 -2636
rect -100 -2717 -84 -2683
rect 84 -2717 100 -2683
rect -100 -2733 100 -2717
<< polycont >>
rect -84 2683 84 2717
rect -84 955 84 989
rect -84 847 84 881
rect -84 -881 84 -847
rect -84 -989 84 -955
rect -84 -2717 84 -2683
<< locali >>
rect -260 2785 -164 2819
rect 164 2785 260 2819
rect -260 2723 -226 2785
rect 226 2723 260 2785
rect -100 2683 -84 2717
rect 84 2683 100 2717
rect -146 2624 -112 2640
rect -146 1032 -112 1048
rect 112 2624 146 2640
rect 112 1032 146 1048
rect -100 955 -84 989
rect 84 955 100 989
rect -100 847 -84 881
rect 84 847 100 881
rect -146 788 -112 804
rect -146 -804 -112 -788
rect 112 788 146 804
rect 112 -804 146 -788
rect -100 -881 -84 -847
rect 84 -881 100 -847
rect -100 -989 -84 -955
rect 84 -989 100 -955
rect -146 -1048 -112 -1032
rect -146 -2640 -112 -2624
rect 112 -1048 146 -1032
rect 112 -2640 146 -2624
rect -100 -2717 -84 -2683
rect 84 -2717 100 -2683
rect -260 -2785 -226 -2723
rect 226 -2785 260 -2723
rect -260 -2819 -164 -2785
rect 164 -2819 260 -2785
<< viali >>
rect -84 2683 84 2717
rect -146 1048 -112 2624
rect 112 1048 146 2624
rect -84 955 84 989
rect -84 847 84 881
rect -146 -788 -112 788
rect 112 -788 146 788
rect -84 -881 84 -847
rect -84 -989 84 -955
rect -146 -2624 -112 -1048
rect 112 -2624 146 -1048
rect -84 -2717 84 -2683
<< metal1 >>
rect -96 2717 96 2723
rect -96 2683 -84 2717
rect 84 2683 96 2717
rect -96 2677 96 2683
rect -152 2624 -106 2636
rect -152 1048 -146 2624
rect -112 1048 -106 2624
rect -152 1036 -106 1048
rect 106 2624 152 2636
rect 106 1048 112 2624
rect 146 1048 152 2624
rect 106 1036 152 1048
rect -96 989 96 995
rect -96 955 -84 989
rect 84 955 96 989
rect -96 949 96 955
rect -96 881 96 887
rect -96 847 -84 881
rect 84 847 96 881
rect -96 841 96 847
rect -152 788 -106 800
rect -152 -788 -146 788
rect -112 -788 -106 788
rect -152 -800 -106 -788
rect 106 788 152 800
rect 106 -788 112 788
rect 146 -788 152 788
rect 106 -800 152 -788
rect -96 -847 96 -841
rect -96 -881 -84 -847
rect 84 -881 96 -847
rect -96 -887 96 -881
rect -96 -955 96 -949
rect -96 -989 -84 -955
rect 84 -989 96 -955
rect -96 -995 96 -989
rect -152 -1048 -106 -1036
rect -152 -2624 -146 -1048
rect -112 -2624 -106 -1048
rect -152 -2636 -106 -2624
rect 106 -1048 152 -1036
rect 106 -2624 112 -1048
rect 146 -2624 152 -1048
rect 106 -2636 152 -2624
rect -96 -2683 96 -2677
rect -96 -2717 -84 -2683
rect 84 -2717 96 -2683
rect -96 -2723 96 -2717
<< properties >>
string FIXED_BBOX -243 -2802 243 2802
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8.0 l 1.0 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
