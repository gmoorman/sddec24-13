magic
tech sky130B
magscale 1 2
timestamp 1734635153
<< nwell >>
rect -216 -1350 4080 1750
<< pwell >>
rect 3700 -1378 3750 -1364
rect -216 -3058 3750 -1378
rect -214 -3068 3750 -3058
<< mvpsubdiff >>
rect -150 -1442 3684 -1430
rect -150 -1542 24 -1442
rect 3510 -1542 3684 -1442
rect -150 -1554 3684 -1542
rect -150 -1604 -26 -1554
rect -150 -2828 -138 -1604
rect -38 -2828 -26 -1604
rect -150 -2878 -26 -2828
rect 3560 -1604 3684 -1554
rect 3560 -2828 3572 -1604
rect 3672 -2828 3684 -1604
rect 3560 -2878 3684 -2828
rect -150 -2890 3684 -2878
rect -150 -2990 24 -2890
rect 3510 -2990 3684 -2890
rect -150 -3002 3684 -2990
<< mvnsubdiff >>
rect -150 1672 4014 1684
rect -150 1572 24 1672
rect 3840 1572 4014 1672
rect -150 1560 4014 1572
rect -150 1510 -26 1560
rect -150 -1104 -138 1510
rect -38 -1104 -26 1510
rect -150 -1154 -26 -1104
rect 3890 1510 4014 1560
rect 3890 -1104 3902 1510
rect 4002 -1104 4014 1510
rect 3890 -1154 4014 -1104
rect -150 -1166 4014 -1154
rect -150 -1266 24 -1166
rect 3840 -1266 4014 -1166
rect -150 -1278 4014 -1266
<< mvpsubdiffcont >>
rect 24 -1542 3510 -1442
rect -138 -2828 -38 -1604
rect 3572 -2828 3672 -1604
rect 24 -2990 3510 -2890
<< mvnsubdiffcont >>
rect 24 1572 3840 1672
rect -138 -1104 -38 1510
rect 3902 -1104 4002 1510
rect 24 -1266 3840 -1166
<< locali >>
rect -138 1510 -38 1672
rect -138 -1266 -38 -1104
rect 3902 1510 4002 1672
rect 3902 -1266 4002 -1104
rect -138 -1604 -38 -1442
rect -138 -2990 -38 -2828
rect 3572 -1604 3672 -1442
rect 3572 -2990 3672 -2828
<< viali >>
rect -38 1572 24 1672
rect 24 1572 3840 1672
rect 3840 1572 3902 1672
rect -138 -1029 -38 1435
rect 3902 -1029 4002 1435
rect -38 -1266 24 -1166
rect 24 -1266 3840 -1166
rect 3840 -1266 3902 -1166
rect -38 -1542 24 -1442
rect 24 -1542 3510 -1442
rect 3510 -1542 3572 -1442
rect -138 -2823 -38 -1609
rect 3572 -2823 3672 -1609
rect -38 -2990 24 -2890
rect 24 -2990 3510 -2890
rect 3510 -2990 3572 -2890
<< metal1 >>
rect -144 1672 4008 1678
rect -144 1572 -38 1672
rect 3902 1572 4008 1672
rect -144 1566 4008 1572
rect -144 1435 -32 1566
rect -144 -1029 -138 1435
rect -38 -1029 -32 1435
rect 568 1266 578 1566
rect 716 1358 768 1368
rect 716 1296 768 1306
rect 724 1142 758 1296
rect 3286 1266 3296 1566
rect 3896 1435 4008 1566
rect 102 1106 3628 1142
rect 310 1004 350 1106
rect 24 936 34 988
rect 86 936 96 988
rect 412 936 422 988
rect 474 936 484 988
rect 664 936 674 988
rect 726 936 736 988
rect 800 936 810 988
rect 862 936 872 988
rect 1052 936 1062 988
rect 1114 936 1124 988
rect 1188 936 1198 988
rect 1250 936 1260 988
rect 1440 936 1450 988
rect 1502 936 1512 988
rect 1576 936 1586 988
rect 1638 936 1648 988
rect 1828 936 1838 988
rect 1890 936 1900 988
rect 1964 936 1974 988
rect 2026 936 2036 988
rect 2216 936 2226 988
rect 2278 936 2288 988
rect 2352 936 2362 988
rect 2414 936 2424 988
rect 2604 936 2614 988
rect 2666 936 2676 988
rect 2740 936 2750 988
rect 2802 936 2812 988
rect 2992 936 3002 988
rect 3054 936 3064 988
rect 3128 936 3138 988
rect 3190 936 3200 988
rect 3380 936 3390 988
rect 3516 936 3526 988
rect 3578 936 3588 988
rect 3532 -110 3566 72
rect 664 -172 674 -120
rect 726 -172 736 -120
rect 1052 -172 1062 -120
rect 1114 -172 1124 -120
rect 1440 -172 1450 -120
rect 1502 -172 1512 -120
rect 1576 -172 1586 -120
rect 1638 -172 1648 -120
rect 1828 -172 1838 -120
rect 1890 -172 1900 -120
rect 2216 -172 2226 -120
rect 2278 -172 2288 -120
rect 2604 -172 2614 -120
rect 2666 -172 2676 -120
rect 2992 -172 3002 -120
rect 3054 -172 3064 -120
rect 3380 -172 3390 -120
rect 412 -362 422 -310
rect 474 -362 484 -310
rect 800 -362 810 -310
rect 862 -362 872 -310
rect 1188 -362 1198 -310
rect 1250 -362 1260 -310
rect 1576 -362 1586 -310
rect 1638 -362 1648 -310
rect 1964 -362 1974 -310
rect 2026 -362 2036 -310
rect 2352 -362 2362 -310
rect 2414 -362 2424 -310
rect 2740 -362 2750 -310
rect 2802 -362 2812 -310
rect 3128 -362 3138 -310
rect 3190 -362 3200 -310
rect -144 -1160 -32 -1029
rect 730 -1080 740 -1068
rect 490 -1114 740 -1080
rect 730 -1120 740 -1114
rect 792 -1080 802 -1068
rect 3058 -1080 3068 -1066
rect 792 -1114 1822 -1080
rect 792 -1120 802 -1114
rect 2042 -1116 3068 -1080
rect 3058 -1118 3068 -1116
rect 3120 -1080 3130 -1066
rect 3120 -1116 3374 -1080
rect 3656 -1114 3700 1142
rect 3768 936 3778 988
rect 3830 936 3840 988
rect 3768 -170 3778 -118
rect 3830 -170 3840 -118
rect 3896 -1029 3902 1435
rect 4002 -1029 4008 1435
rect 3120 -1118 3130 -1116
rect 3896 -1160 4008 -1029
rect -144 -1166 4008 -1160
rect -144 -1266 -38 -1166
rect 3902 -1266 4008 -1166
rect -144 -1272 4008 -1266
rect -144 -1442 3678 -1436
rect -144 -1542 -38 -1442
rect 3572 -1542 3678 -1442
rect -144 -1548 3678 -1542
rect -144 -1609 -32 -1548
rect -144 -2823 -138 -1609
rect -38 -2823 -32 -1609
rect 412 -1614 1648 -1586
rect 412 -1666 422 -1614
rect 474 -1666 484 -1614
rect 800 -1666 810 -1614
rect 862 -1666 872 -1614
rect 1190 -1666 1200 -1614
rect 1252 -1666 1262 -1614
rect 1576 -1666 1586 -1614
rect 1638 -1666 1648 -1614
rect 1966 -1614 3198 -1586
rect 1966 -1666 1976 -1614
rect 2028 -1666 2038 -1614
rect 2352 -1666 2362 -1614
rect 2414 -1666 2424 -1614
rect 2740 -1666 2750 -1614
rect 2802 -1666 2812 -1614
rect 3126 -1666 3136 -1614
rect 3188 -1666 3198 -1614
rect 3566 -1609 3678 -1548
rect 664 -2084 674 -2032
rect 726 -2084 736 -2032
rect 1052 -2084 1062 -2032
rect 1114 -2084 1124 -2032
rect 1442 -2084 1452 -2032
rect 1504 -2084 1514 -2032
rect 1828 -2084 1838 -2032
rect 1890 -2084 1900 -2032
rect 2218 -2084 2228 -2032
rect 2280 -2084 2290 -2032
rect 2604 -2084 2614 -2032
rect 2666 -2084 2676 -2032
rect 2992 -2084 3002 -2032
rect 3054 -2084 3064 -2032
rect 3378 -2084 3388 -2032
rect 3440 -2084 3450 -2032
rect 446 -2492 480 -2430
rect 2000 -2492 2034 -2428
rect 446 -2526 1780 -2492
rect 2000 -2526 3334 -2492
rect -144 -2884 -32 -2823
rect 568 -2884 578 -2584
rect 2956 -2884 2966 -2584
rect 3566 -2823 3572 -1609
rect 3672 -2823 3678 -1609
rect 3566 -2884 3678 -2823
rect -144 -2890 3678 -2884
rect -144 -2990 -38 -2890
rect 3572 -2990 3678 -2890
rect -144 -2996 3678 -2990
<< via1 >>
rect -32 1266 568 1566
rect 716 1306 768 1358
rect 3296 1266 3896 1566
rect 34 936 86 988
rect 422 936 474 988
rect 674 936 726 988
rect 810 936 862 988
rect 1062 936 1114 988
rect 1198 936 1250 988
rect 1450 936 1502 988
rect 1586 936 1638 988
rect 1838 936 1890 988
rect 1974 936 2026 988
rect 2226 936 2278 988
rect 2362 936 2414 988
rect 2614 936 2666 988
rect 2750 936 2802 988
rect 3002 936 3054 988
rect 3138 936 3190 988
rect 3390 936 3442 988
rect 3526 936 3578 988
rect 674 -172 726 -120
rect 1062 -172 1114 -120
rect 1450 -172 1502 -120
rect 1586 -172 1638 -120
rect 1838 -172 1890 -120
rect 2226 -172 2278 -120
rect 2614 -172 2666 -120
rect 3002 -172 3054 -120
rect 3390 -172 3442 -120
rect 422 -362 474 -310
rect 810 -362 862 -310
rect 1198 -362 1250 -310
rect 1586 -362 1638 -310
rect 1974 -362 2026 -310
rect 2362 -362 2414 -310
rect 2750 -362 2802 -310
rect 3138 -362 3190 -310
rect 740 -1120 792 -1068
rect 3068 -1118 3120 -1066
rect 3778 936 3830 988
rect 3778 -170 3830 -118
rect 422 -1666 474 -1614
rect 810 -1666 862 -1614
rect 1200 -1666 1252 -1614
rect 1586 -1666 1638 -1614
rect 1976 -1666 2028 -1614
rect 2362 -1666 2414 -1614
rect 2750 -1666 2802 -1614
rect 3136 -1666 3188 -1614
rect 674 -2084 726 -2032
rect 1062 -2084 1114 -2032
rect 1452 -2084 1504 -2032
rect 1838 -2084 1890 -2032
rect 2228 -2084 2280 -2032
rect 2614 -2084 2666 -2032
rect 3002 -2084 3054 -2032
rect 3388 -2084 3440 -2032
rect -32 -2884 568 -2584
rect 2966 -2884 3566 -2584
<< metal2 >>
rect -32 1566 568 1576
rect 3296 1566 3896 1576
rect 778 1358 838 1364
rect 706 1306 716 1358
rect 768 1306 838 1358
rect 778 1304 838 1306
rect -32 1256 568 1266
rect 3296 1256 3896 1266
rect 40 1152 74 1256
rect 204 1254 238 1256
rect 40 1122 3566 1152
rect 40 998 74 1122
rect 428 998 462 1122
rect 816 998 850 1122
rect 1204 998 1238 1122
rect 1592 998 1626 1122
rect 1980 998 2014 1122
rect 2368 998 2402 1122
rect 2756 998 2790 1122
rect 3144 998 3178 1122
rect 3532 998 3566 1122
rect 34 988 86 998
rect 34 926 86 936
rect 422 988 474 998
rect 422 926 474 936
rect 674 988 726 998
rect 674 926 726 936
rect 810 988 862 998
rect 810 926 862 936
rect 1062 988 1114 998
rect 1062 926 1114 936
rect 1198 988 1250 998
rect 1198 926 1250 936
rect 1450 988 1502 998
rect 1450 926 1502 936
rect 1586 988 1638 998
rect 1586 926 1638 936
rect 1838 988 1890 998
rect 1838 926 1890 936
rect 1974 988 2026 998
rect 1974 926 2026 936
rect 2226 988 2278 998
rect 2226 926 2278 936
rect 2362 988 2414 998
rect 2362 926 2414 936
rect 2614 988 2666 998
rect 2614 926 2666 936
rect 2750 988 2802 998
rect 2750 926 2802 936
rect 3002 988 3054 998
rect 3002 926 3054 936
rect 3138 988 3190 998
rect 3138 926 3190 936
rect 3390 988 3442 998
rect 3390 926 3442 936
rect 3526 988 3578 998
rect 3526 926 3578 936
rect 3778 988 3830 998
rect 3778 926 3830 936
rect 686 28 720 926
rect 1074 28 1108 926
rect 1462 28 1496 926
rect 1850 28 1884 926
rect 2238 28 2272 926
rect 2626 28 2660 926
rect 3014 28 3048 926
rect 3402 28 3436 926
rect 3790 28 3824 926
rect 686 0 3824 28
rect 686 -110 720 0
rect 1074 -110 1108 0
rect 1462 -110 1496 0
rect 1850 -110 1884 0
rect 2238 -110 2272 0
rect 2626 -110 2660 0
rect 3014 -110 3048 0
rect 3402 -110 3436 0
rect 3790 -108 3824 0
rect 674 -120 726 -110
rect 674 -182 726 -172
rect 1062 -120 1114 -110
rect 1062 -182 1114 -172
rect 1450 -120 1502 -110
rect 1450 -178 1502 -172
rect 1586 -120 1638 -110
rect 1586 -182 1638 -172
rect 1838 -120 1890 -110
rect 1838 -182 1890 -172
rect 2226 -120 2278 -110
rect 2226 -182 2278 -172
rect 2614 -120 2666 -110
rect 2614 -178 2666 -172
rect 3002 -120 3054 -110
rect 3002 -182 3054 -172
rect 3390 -120 3442 -110
rect 3390 -182 3442 -172
rect 3778 -118 3830 -108
rect 3778 -180 3830 -170
rect 422 -310 474 -300
rect 810 -310 862 -300
rect 1198 -310 1250 -300
rect 1586 -310 1638 -300
rect 474 -362 810 -310
rect 862 -362 1198 -310
rect 1250 -362 1586 -310
rect 422 -372 474 -362
rect 810 -372 862 -362
rect 1198 -372 1250 -362
rect 1586 -372 1638 -362
rect 1974 -310 2026 -300
rect 2362 -310 2414 -300
rect 2750 -310 2802 -300
rect 3138 -310 3190 -300
rect 2026 -362 2362 -310
rect 2414 -362 2750 -310
rect 2802 -362 3138 -310
rect 1974 -372 2026 -362
rect 2362 -372 2414 -362
rect 2750 -372 2802 -362
rect 3138 -372 3190 -362
rect 740 -1068 792 -1058
rect 740 -1130 792 -1120
rect 736 -1190 796 -1130
rect 1208 -1338 1242 -372
rect 2368 -1338 2402 -372
rect 3068 -1066 3120 -1056
rect 3068 -1128 3120 -1118
rect 3064 -1188 3124 -1128
rect 1194 -1398 1254 -1338
rect 2356 -1398 2416 -1338
rect 1208 -1604 1242 -1398
rect 422 -1614 474 -1604
rect 422 -1676 474 -1666
rect 810 -1614 862 -1604
rect 810 -1676 862 -1666
rect 1200 -1614 1252 -1604
rect 1200 -1676 1252 -1666
rect 1586 -1614 1638 -1604
rect 1586 -1676 1638 -1666
rect 1976 -1614 2028 -1604
rect 2368 -1608 2402 -1398
rect 1976 -1676 2028 -1666
rect 2362 -1614 2414 -1608
rect 2362 -1676 2414 -1666
rect 2750 -1614 2802 -1604
rect 2750 -1676 2802 -1666
rect 3136 -1614 3188 -1604
rect 3136 -1676 3188 -1666
rect 822 -1790 856 -1676
rect 674 -2032 726 -2022
rect 1062 -2032 1114 -2022
rect 726 -2074 1062 -2040
rect 674 -2094 726 -2084
rect 1452 -2032 1504 -2022
rect 1114 -2074 1452 -2040
rect 1062 -2094 1114 -2084
rect 1838 -2032 1890 -2022
rect 1504 -2074 1838 -2040
rect 1452 -2094 1504 -2084
rect 2228 -2032 2280 -2022
rect 1890 -2074 2228 -2040
rect 1838 -2094 1890 -2084
rect 2614 -2032 2666 -2022
rect 2280 -2074 2614 -2040
rect 2228 -2094 2280 -2084
rect 3002 -2032 3054 -2022
rect 2666 -2074 3002 -2040
rect 2614 -2094 2666 -2084
rect 3388 -2032 3440 -2022
rect 3054 -2074 3388 -2040
rect 3002 -2094 3054 -2084
rect 3388 -2094 3440 -2084
rect -32 -2584 568 -2574
rect 686 -2598 720 -2094
rect 568 -2628 720 -2598
rect 2966 -2584 3566 -2574
rect -32 -2894 568 -2884
rect 2966 -2894 3566 -2884
<< via2 >>
rect -32 1266 568 1566
rect 3296 1266 3896 1566
rect -32 -2884 568 -2584
rect 2966 -2884 3566 -2584
<< metal3 >>
rect -42 1566 578 1571
rect -42 1266 -32 1566
rect 568 1266 578 1566
rect -42 1261 578 1266
rect 3286 1566 3906 1571
rect 3286 1266 3296 1566
rect 3896 1266 3906 1566
rect 3286 1261 3906 1266
rect -42 -2584 578 -2579
rect -42 -2884 -32 -2584
rect 568 -2884 578 -2584
rect -42 -2889 578 -2884
rect 2956 -2584 3576 -2579
rect 2956 -2884 2966 -2584
rect 3566 -2884 3576 -2584
rect 2956 -2889 3576 -2884
<< via3 >>
rect -32 1266 568 1566
rect 3296 1266 3896 1566
rect -32 -2884 568 -2584
rect 2966 -2884 3566 -2584
<< metal4 >>
rect -33 1566 569 1567
rect -33 1266 -32 1566
rect 568 1266 569 1566
rect -33 1265 569 1266
rect 3295 1566 3897 1567
rect 3295 1266 3296 1566
rect 3896 1266 3897 1566
rect 3295 1265 3897 1266
rect -33 -2584 569 -2583
rect -33 -2884 -32 -2584
rect 568 -2884 569 -2584
rect -33 -2885 569 -2884
rect 2965 -2584 3567 -2583
rect 2965 -2884 2966 -2584
rect 3566 -2884 3567 -2584
rect 2965 -2885 3567 -2884
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_0 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold/gds_isolate
timestamp 1734209266
transform 1 0 2902 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_1
timestamp 1734209266
transform 1 0 574 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_2
timestamp 1734209266
transform 1 0 962 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_3
timestamp 1734209266
transform 1 0 1352 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_4
timestamp 1734209266
transform 1 0 1738 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_5
timestamp 1734209266
transform 1 0 2128 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_6
timestamp 1734209266
transform 1 0 2514 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_GKZ9Z2  sky130_fd_pr__nfet_01v8_GKZ9Z2_7
timestamp 1734209266
transform 1 0 3288 0 1 -2085
box -158 -457 158 457
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_0 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold/gds_isolate
timestamp 1734634369
transform 1 0 574 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_1
timestamp 1734634369
transform 1 0 962 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_2
timestamp 1734634369
transform 1 0 1350 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_3
timestamp 1734634369
transform 1 0 1738 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_4
timestamp 1734634369
transform 1 0 2126 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_5
timestamp 1734634369
transform 1 0 2514 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_6
timestamp 1734634369
transform 1 0 2902 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_7
timestamp 1734634369
transform 1 0 3290 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_8
timestamp 1734634369
transform 1 0 3678 0 1 -570
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_0 ~/caravel_pls_man_analog/caravel_user_project_analog/mag/comparator_hold/gds_isolate
timestamp 1734634369
transform 1 0 3678 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_1
timestamp 1734634369
transform 1 0 962 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_2
timestamp 1734634369
transform 1 0 186 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_3
timestamp 1734634369
transform 1 0 1350 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_4
timestamp 1734634369
transform 1 0 1738 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_5
timestamp 1734634369
transform 1 0 2126 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_6
timestamp 1734634369
transform 1 0 2514 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_7
timestamp 1734634369
transform 1 0 2902 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_8
timestamp 1734634369
transform 1 0 3290 0 1 596
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_9
timestamp 1734634369
transform 1 0 574 0 1 596
box -194 -598 194 564
<< labels >>
rlabel metal2 778 1304 838 1364 1 curr_in
port 3 n
rlabel metal2 3064 -1188 3124 -1128 1 Vinplus
port 5 n
rlabel metal2 1194 -1398 1254 -1338 1 Viominus
port 6 n
rlabel metal2 2356 -1398 2416 -1338 1 Vioplus
port 7 n
rlabel metal2 736 -1190 796 -1130 1 Vinminus
port 8 n
rlabel via2 198 -2774 258 -2714 1 VSS
port 1 n
rlabel via2 194 1338 254 1398 1 VDD
port 2 n
<< properties >>
string FIXED_BBOX -302 -2932 3572 -1484
<< end >>
