magic
tech sky130B
magscale 1 2
timestamp 1733716281
<< nwell >>
rect -1116 9486 37204 9588
rect -1526 9356 -728 9438
<< pwell >>
rect 13156 50 13186 6572
rect 26314 50 26344 6572
rect -4388 -718 -4358 -76
rect -1486 -376 -1446 -44
rect -454 -52 37866 50
rect -2 -718 28 -76
rect 2900 -398 2940 -52
rect 7286 -398 7326 -52
rect 11672 -398 11712 -52
rect 13156 -718 13186 -52
rect 16058 -398 16098 -52
rect 20444 -398 20484 -52
rect 24830 -398 24870 -52
rect 26314 -718 26344 -52
rect 29216 -398 29256 -52
rect 33602 -398 33642 -52
rect 37988 -398 38028 -44
rect 39472 -718 39502 6572
rect 42374 -398 42414 -44
rect 46760 -398 46800 -44
rect 51146 -400 51186 -46
rect 52630 -720 52660 6570
rect 61550 2214 61620 2268
rect 55532 -400 55572 -46
rect 59942 -400 59982 -46
rect 64300 -402 64340 -48
<< metal1 >>
rect -1116 9486 65598 9588
rect -454 -44 42390 50
rect 46776 -44 65598 50
rect -1486 -376 -1446 -44
rect -454 -52 42414 -44
rect 2900 -398 2940 -52
rect 7286 -398 7326 -52
rect 11672 -398 11712 -52
rect 16058 -398 16098 -52
rect 20444 -398 20484 -52
rect 24830 -398 24870 -52
rect 29216 -398 29256 -52
rect 33602 -398 33642 -52
rect 37988 -398 38028 -52
rect 42374 -398 42414 -52
rect 46760 -52 65598 -44
rect 46760 -398 46800 -52
rect 51146 -400 51186 -52
rect 55532 -400 55572 -52
rect 59942 -400 59982 -52
rect 64300 -402 64340 -52
<< metal2 >>
rect -1264 9854 -1254 9926
rect -1182 9854 -1172 9926
rect 3122 9854 3132 9926
rect 3204 9854 3214 9926
rect 7508 9856 7518 9928
rect 7590 9856 7600 9928
rect 11894 9856 11904 9928
rect 11976 9856 11986 9928
rect 16280 9852 16290 9924
rect 16362 9852 16372 9924
rect 20668 9868 20678 9940
rect 20750 9868 20760 9940
rect 25052 9856 25062 9928
rect 25134 9856 25144 9928
rect 35926 9926 38290 9928
rect 29438 9852 29448 9924
rect 29520 9852 29530 9924
rect 34222 9906 34232 9922
rect 33888 9850 34232 9906
rect 34304 9850 34314 9922
rect 35834 9854 35844 9926
rect 35916 9856 38290 9926
rect 35916 9854 35926 9856
rect 40286 9848 40296 9920
rect 40368 9848 42692 9920
rect 46980 9854 46990 9926
rect 47062 9854 47072 9926
rect 51368 9856 51378 9928
rect 51450 9856 51460 9928
rect 55754 9850 55764 9922
rect 55836 9850 55846 9922
rect 60142 9850 60152 9922
rect 60224 9850 60234 9922
rect 64526 9850 64536 9922
rect 64608 9850 64618 9922
rect -1032 6660 -960 6670
rect -1032 6578 -960 6588
rect 3354 6662 3426 6672
rect 3354 6580 3426 6590
rect 7744 6662 7816 6672
rect 7744 6580 7816 6590
rect 12130 6662 12202 6672
rect 12130 6580 12202 6590
rect 16514 6658 16586 6668
rect 16514 6576 16586 6586
rect 20900 6662 20972 6672
rect 20900 6580 20972 6590
rect 25284 6660 25356 6670
rect 25284 6578 25356 6588
rect 29672 6662 29744 6672
rect 29672 6580 29744 6590
rect 34058 6660 34130 6670
rect 34058 6578 34130 6588
rect 38444 6662 38516 6672
rect 38444 6580 38516 6590
rect 42830 6660 42902 6670
rect 42830 6578 42902 6588
rect 47216 6658 47288 6668
rect 47216 6576 47288 6586
rect 51602 6660 51674 6670
rect 51602 6578 51674 6588
rect 55988 6662 56060 6672
rect 55988 6580 56060 6590
rect 60372 6658 60444 6668
rect 60372 6576 60444 6586
rect 64760 6658 64832 6668
rect 64760 6576 64832 6586
rect -4438 2218 -4140 2272
rect -52 2218 246 2272
rect 4334 2218 4632 2272
rect 8720 2218 9018 2272
rect 13106 2218 13332 2272
rect 17492 2218 17790 2272
rect 21878 2218 22176 2272
rect 26264 2218 26490 2272
rect 30650 2218 30948 2272
rect 35036 2218 35334 2272
rect 39422 2218 39648 2272
rect 43808 2218 44106 2272
rect -4438 -108 -4358 2218
rect -524 2116 -246 2166
rect -4388 -682 -4358 -108
rect -284 -682 -246 2116
rect -52 -108 28 2218
rect 3862 2116 4140 2166
rect -4388 -718 -3160 -682
rect -3052 -718 -246 -682
rect -2 -682 28 -108
rect 4102 -682 4140 2116
rect 4334 -108 4414 2218
rect 8248 2116 8526 2166
rect -2 -718 1226 -682
rect 1334 -718 4140 -682
rect 4384 -682 4414 -108
rect 8488 -682 8526 2116
rect 8720 -108 8800 2218
rect 12634 2116 12912 2166
rect 4384 -718 5612 -682
rect 5720 -718 8526 -682
rect 8770 -682 8800 -108
rect 12874 -682 12912 2116
rect 13106 -108 13186 2218
rect 17064 2116 17298 2166
rect 8770 -718 9998 -682
rect 10106 -718 12912 -682
rect 13156 -682 13186 -108
rect 17260 -682 17298 2116
rect 17492 -108 17572 2218
rect 21406 2116 21684 2166
rect 13156 -718 14384 -682
rect 14492 -718 17298 -682
rect 17542 -682 17572 -108
rect 21646 -682 21684 2116
rect 21878 -108 21958 2218
rect 25792 2116 26070 2166
rect 17542 -718 18770 -682
rect 18878 -718 21684 -682
rect 21928 -682 21958 -108
rect 26032 -682 26070 2116
rect 26264 -108 26344 2218
rect 30222 2116 30456 2166
rect 21928 -718 23156 -682
rect 23264 -718 26070 -682
rect 26314 -682 26344 -108
rect 30418 -682 30456 2116
rect 30650 -108 30730 2218
rect 34564 2116 34842 2166
rect 26314 -718 27542 -682
rect 27650 -718 30456 -682
rect 30700 -682 30730 -108
rect 34804 -682 34842 2116
rect 35036 -108 35116 2218
rect 38950 2116 39228 2166
rect 30700 -718 31928 -682
rect 32036 -718 34842 -682
rect 35086 -682 35116 -108
rect 39190 -682 39228 2116
rect 39422 -108 39502 2218
rect 43380 2116 43614 2166
rect 35086 -718 36314 -682
rect 36422 -718 39228 -682
rect 39472 -682 39502 -108
rect 43576 -682 43614 2116
rect 43808 -108 43888 2218
rect 48194 2216 48492 2270
rect 52580 2216 52806 2270
rect 56966 2216 57264 2270
rect 47722 2116 48000 2166
rect 39472 -718 40700 -682
rect 40808 -718 43614 -682
rect 43858 -682 43888 -108
rect 47962 -682 48000 2116
rect 48194 -110 48274 2216
rect 52108 2114 52386 2164
rect 43858 -718 45086 -682
rect 45194 -718 48000 -682
rect 48244 -684 48274 -110
rect 52348 -684 52386 2114
rect 52580 -110 52660 2216
rect 56538 2114 56772 2164
rect 48244 -720 49472 -684
rect 49580 -720 52386 -684
rect 52630 -684 52660 -110
rect 56734 -684 56772 2114
rect 56966 -110 57046 2216
rect 61324 2214 61620 2268
rect 60880 2114 61158 2164
rect 52630 -720 53858 -684
rect 53966 -720 56772 -684
rect 57016 -684 57046 -110
rect 61120 -684 61158 2114
rect 61324 -112 61404 2214
rect 64648 2092 64676 2144
rect 65282 2112 65516 2162
rect 57016 -720 58244 -684
rect 58352 -720 61158 -684
rect 61374 -686 61404 -112
rect 65478 -686 65516 2112
rect 61374 -722 62602 -686
rect 62710 -722 65516 -686
<< via2 >>
rect -1254 9854 -1182 9926
rect 3132 9854 3204 9926
rect 7518 9856 7590 9928
rect 11904 9856 11976 9928
rect 16290 9852 16362 9924
rect 20678 9868 20750 9940
rect 25062 9856 25134 9928
rect 29448 9852 29520 9924
rect 34232 9850 34304 9922
rect 35844 9854 35916 9926
rect 40296 9848 40368 9920
rect 46990 9854 47062 9926
rect 51378 9856 51450 9928
rect 55764 9850 55836 9922
rect 60152 9850 60224 9922
rect 64536 9850 64608 9922
rect -1032 6588 -960 6660
rect 3354 6590 3426 6662
rect 7744 6590 7816 6662
rect 12130 6590 12202 6662
rect 16514 6586 16586 6658
rect 20900 6590 20972 6662
rect 25284 6588 25356 6660
rect 29672 6590 29744 6662
rect 34058 6588 34130 6660
rect 38444 6590 38516 6662
rect 42830 6588 42902 6660
rect 47216 6586 47288 6658
rect 51602 6588 51674 6660
rect 55988 6590 56060 6662
rect 60372 6586 60444 6658
rect 64760 6586 64832 6658
<< metal3 >>
rect 32996 11810 33028 11928
rect 32996 10904 33058 11810
rect 33784 11594 33820 11714
rect -1254 10844 33058 10904
rect -1254 9936 -1180 10844
rect 33210 10784 33272 11108
rect 3118 10724 33272 10784
rect 3132 9936 3204 10724
rect 33482 10664 33544 11110
rect 7504 10604 33544 10664
rect 7518 9938 7590 10604
rect 33754 10542 33820 11594
rect 11892 10482 33820 10542
rect 11904 9938 11976 10482
rect 34026 10422 34092 11108
rect 16276 10362 34094 10422
rect -1259 9926 -1177 9936
rect -1259 9854 -1254 9926
rect -1182 9854 -1177 9926
rect -1259 9844 -1177 9854
rect 3127 9926 3209 9936
rect 3127 9854 3132 9926
rect 3204 9854 3209 9926
rect 3127 9844 3209 9854
rect 7513 9928 7595 9938
rect 7513 9856 7518 9928
rect 7590 9856 7595 9928
rect 7513 9846 7595 9856
rect 11899 9928 11981 9938
rect 16290 9934 16362 10362
rect 20678 10300 34112 10302
rect 34294 10300 34360 11116
rect 20678 10238 34360 10300
rect 20678 9950 20750 10238
rect 34570 10178 34636 11116
rect 25042 10118 34636 10178
rect 20673 9940 20755 9950
rect 11899 9856 11904 9928
rect 11976 9856 11981 9928
rect 11899 9846 11981 9856
rect 16285 9924 16367 9934
rect 16285 9852 16290 9924
rect 16362 9852 16367 9924
rect 20673 9868 20678 9940
rect 20750 9868 20755 9940
rect 25062 9938 25142 10118
rect 34840 10058 34906 11116
rect 29434 9998 34906 10058
rect 35110 10874 35176 11110
rect 35430 10878 35496 11116
rect 35700 10878 35766 11118
rect 35980 10880 36046 11110
rect 36252 10882 36318 11110
rect 36524 10882 36590 11110
rect 29434 9994 34640 9998
rect 20673 9858 20755 9868
rect 25057 9928 25142 9938
rect 16285 9842 16367 9852
rect 25057 9856 25062 9928
rect 25134 9858 25142 9928
rect 29442 9924 29526 9994
rect 25134 9856 25139 9858
rect 25057 9846 25139 9856
rect 29442 9854 29448 9924
rect 29443 9852 29448 9854
rect 29520 9854 29526 9924
rect 34227 9922 34309 9932
rect 29520 9852 29525 9854
rect 29443 9842 29525 9852
rect 34227 9850 34232 9922
rect 34304 9850 34309 9922
rect 34227 9840 34309 9850
rect 34230 9780 34308 9840
rect 34230 9778 34958 9780
rect 35110 9778 35178 10874
rect 35430 9784 35506 10878
rect 35700 10056 35776 10878
rect 35980 10176 36050 10880
rect 36252 10302 36322 10882
rect 36524 10424 36594 10882
rect 36796 10546 36866 11062
rect 37072 10670 37142 11068
rect 37072 10668 37898 10670
rect 37072 10608 64640 10668
rect 36796 10544 37622 10546
rect 36796 10484 60236 10544
rect 36524 10422 37350 10424
rect 36524 10362 55836 10422
rect 36252 10296 37058 10302
rect 36252 10236 51460 10296
rect 51062 10234 51460 10236
rect 35980 10116 47074 10176
rect 35700 9996 40368 10056
rect 35839 9926 35921 9936
rect 40296 9930 40368 9996
rect 46990 9936 47060 10116
rect 51376 9938 51460 10234
rect 35839 9854 35844 9926
rect 35916 9854 35921 9926
rect 35839 9844 35921 9854
rect 40291 9920 40373 9930
rect 40291 9848 40296 9920
rect 40368 9848 40373 9920
rect 35842 9784 35916 9844
rect 40291 9838 40373 9848
rect 46985 9926 47067 9936
rect 46985 9854 46990 9926
rect 47062 9854 47067 9926
rect 46985 9844 47067 9854
rect 51373 9928 51460 9938
rect 55764 9932 55836 10362
rect 60152 9932 60236 10484
rect 64536 9932 64612 10608
rect 51373 9856 51378 9928
rect 51450 9856 51460 9928
rect 55759 9922 55841 9932
rect 51373 9846 51455 9856
rect 55759 9850 55764 9922
rect 55836 9850 55841 9922
rect 55759 9840 55841 9850
rect 60147 9922 60236 9932
rect 60147 9850 60152 9922
rect 60224 9850 60236 9922
rect 64531 9922 64613 9932
rect 64531 9850 64536 9922
rect 64608 9850 64613 9922
rect 60147 9840 60229 9850
rect 64531 9840 64613 9850
rect 34230 9718 35176 9778
rect 35430 9720 35920 9784
rect -1042 6660 -950 6665
rect 3344 6662 3436 6667
rect -1042 6658 -1032 6660
rect -4742 6588 -1032 6658
rect -960 6658 -898 6660
rect 3344 6658 3354 6662
rect -960 6590 3354 6658
rect 3426 6658 3436 6662
rect 7734 6662 7826 6667
rect 7734 6658 7744 6662
rect 3426 6590 7744 6658
rect 7816 6658 7826 6662
rect 12120 6662 12212 6667
rect 12120 6658 12130 6662
rect 7816 6590 12130 6658
rect 12202 6658 12212 6662
rect 16504 6658 16596 6663
rect 20890 6662 20982 6667
rect 20890 6658 20900 6662
rect 12202 6590 16514 6658
rect -960 6588 16514 6590
rect -4742 6586 16514 6588
rect 16586 6590 20900 6658
rect 20972 6658 20982 6662
rect 25274 6660 25366 6665
rect 25274 6658 25284 6660
rect 20972 6590 25284 6658
rect 16586 6588 25284 6590
rect 25356 6658 25366 6660
rect 29662 6662 29754 6667
rect 29662 6658 29672 6662
rect 25356 6590 29672 6658
rect 29744 6658 29754 6662
rect 34048 6660 34140 6665
rect 34048 6658 34058 6660
rect 29744 6590 34058 6658
rect 25356 6588 34058 6590
rect 34130 6658 34140 6660
rect 38434 6662 38526 6667
rect 38434 6658 38444 6662
rect 34130 6590 38444 6658
rect 38516 6658 38526 6662
rect 42820 6660 42912 6665
rect 42820 6658 42830 6660
rect 38516 6590 42830 6658
rect 34130 6588 42830 6590
rect 42902 6658 42912 6660
rect 47206 6658 47298 6663
rect 51592 6660 51684 6665
rect 51592 6658 51602 6660
rect 42902 6588 47216 6658
rect 16586 6586 47216 6588
rect 47288 6588 51602 6658
rect 51674 6658 51684 6660
rect 55978 6662 56070 6667
rect 55978 6658 55988 6662
rect 51674 6590 55988 6658
rect 56060 6658 56070 6662
rect 60362 6658 60454 6663
rect 64750 6658 64842 6663
rect 56060 6590 60372 6658
rect 51674 6588 60372 6590
rect 47288 6586 60372 6588
rect 60444 6586 64760 6658
rect 64832 6586 64842 6658
rect -1042 6583 -950 6586
rect 3344 6585 3436 6586
rect 7734 6585 7826 6586
rect 12120 6585 12212 6586
rect 16504 6581 16596 6586
rect 20890 6585 20982 6586
rect 25274 6583 25366 6586
rect 29662 6585 29754 6586
rect 34048 6583 34140 6586
rect 38434 6585 38526 6586
rect 42820 6583 42912 6586
rect 47206 6581 47298 6586
rect 51592 6583 51684 6586
rect 55978 6585 56070 6586
rect 60362 6581 60454 6586
rect 64750 6581 64842 6586
<< metal4 >>
rect -1528 9356 -728 9438
rect -1528 -1150 -1430 9356
rect -1528 -1240 64412 -1150
use combination_test_DUMMY  combination_test_DUMMY_0
timestamp 1733627311
transform 1 0 53078 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_1
timestamp 1733627311
transform 1 0 446 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_2
timestamp 1733627311
transform 1 0 39920 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_3
timestamp 1733627311
transform 1 0 48692 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_4
timestamp 1733627311
transform 1 0 44306 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_5
timestamp 1733627311
transform 1 0 17990 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_6
timestamp 1733627311
transform 1 0 13604 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_7
timestamp 1733627311
transform 1 0 9218 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_8
timestamp 1733627311
transform 1 0 4832 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_9
timestamp 1733627311
transform 1 0 22376 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_10
timestamp 1733627311
transform 1 0 26762 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_11
timestamp 1733627311
transform 1 0 31148 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_12
timestamp 1733627311
transform 1 0 35534 0 1 8472
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_13
timestamp 1733627311
transform 1 0 57464 0 1 8470
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_14
timestamp 1733627311
transform 1 0 61850 0 1 8470
box -574 -8600 3812 1466
use combination_test_DUMMY  combination_test_DUMMY_15
timestamp 1733627311
transform 1 0 -3940 0 1 8472
box -574 -8600 3812 1466
use Preamp_noBias  Preamp_noBias_0
timestamp 1733704917
transform 0 1 40876 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_1
timestamp 1733704917
transform 0 1 32104 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_2
timestamp 1733704917
transform 0 1 23332 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_3
timestamp 1733704917
transform 0 1 5788 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_4
timestamp 1733704917
transform 0 1 1402 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_5
timestamp 1733704917
transform 0 1 -2984 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_6
timestamp 1733704917
transform 0 1 10174 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_7
timestamp 1733704917
transform 0 1 14560 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_8
timestamp 1733704917
transform 0 1 18946 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_9
timestamp 1733704917
transform 0 1 36490 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_10
timestamp 1733704917
transform 0 1 27718 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_11
timestamp 1733704917
transform 0 1 62802 1 0 -4808
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_12
timestamp 1733704917
transform 0 1 49648 1 0 -4806
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_13
timestamp 1733704917
transform 0 1 54034 1 0 -4806
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_14
timestamp 1733704917
transform 0 1 45262 1 0 -4804
box -240 -1530 4730 1840
use Preamp_noBias  Preamp_noBias_15
timestamp 1733704917
transform 0 1 58444 1 0 -4806
box -240 -1530 4730 1840
use Priority_Encoder_16t4  Priority_Encoder_16t4_0
timestamp 1733649010
transform 0 -1 39050 -1 0 19008
box 0 1812 8000 6112
<< end >>
