magic
tech sky130B
timestamp 1731450402
<< checkpaint >>
rect -630 -1230 730 730
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 TE
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 BE
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 Tfilament_0=3.3e-9
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 area_ox=0.1024e-12
port 3 nsew
<< end >>
