magic
tech sky130B
magscale 1 2
timestamp 1733079491
<< nwell >>
rect -574 -1780 3812 1200
<< pwell >>
rect -574 -8672 3812 -1900
<< nmos >>
rect 264 -3009 294 -2609
rect 544 -3009 574 -2609
rect 824 -3009 854 -2609
rect 1104 -3009 1134 -2609
rect 1384 -3009 1414 -2609
rect 1664 -3009 1694 -2609
rect 1944 -3009 1974 -2609
rect 2224 -3009 2254 -2609
rect 2504 -3009 2534 -2609
rect 2784 -3009 2814 -2609
rect 264 -3829 294 -3429
rect 544 -3829 574 -3429
rect 824 -3829 854 -3429
rect 1104 -3829 1134 -3429
rect 1384 -3829 1414 -3429
rect 1664 -3829 1694 -3429
rect 1944 -3829 1974 -3429
rect 2224 -3829 2254 -3429
rect 2504 -3829 2534 -3429
rect 2784 -3829 2814 -3429
rect 1384 -5109 1414 -4709
rect 1664 -5109 1694 -4709
rect 1383 -5967 1413 -5567
rect 1663 -5967 1693 -5567
rect 264 -6912 294 -6512
rect 544 -6912 574 -6512
rect 824 -6912 854 -6512
rect 1104 -6912 1134 -6512
rect 1384 -6912 1414 -6512
rect 1664 -6912 1694 -6512
rect 1944 -6912 1974 -6512
rect 2224 -6912 2254 -6512
rect 2504 -6912 2534 -6512
rect 2784 -6912 2814 -6512
rect 264 -7610 294 -7210
rect 544 -7610 574 -7210
rect 824 -7610 854 -7210
rect 1104 -7610 1134 -7210
rect 1384 -7610 1414 -7210
rect 1664 -7610 1694 -7210
rect 1944 -7610 1974 -7210
rect 2224 -7610 2254 -7210
rect 2504 -7610 2534 -7210
rect 2784 -7610 2814 -7210
<< pmos >>
rect -15 -200 15 200
rect 265 -200 295 200
rect 545 -200 575 200
rect 825 -200 855 200
rect 1105 -200 1135 200
rect 1385 -200 1415 200
rect 1665 -200 1695 200
rect 1945 -200 1975 200
rect 2225 -200 2255 200
rect 2505 -200 2535 200
rect 2785 -200 2815 200
rect 3065 -200 3095 200
rect -15 -916 15 -516
rect 265 -916 295 -516
rect 545 -916 575 -516
rect 825 -916 855 -516
rect 1105 -916 1135 -516
rect 1385 -916 1415 -516
rect 1665 -916 1695 -516
rect 1945 -916 1975 -516
rect 2225 -916 2255 -516
rect 2505 -916 2535 -516
rect 2785 -916 2815 -516
rect 3065 -916 3095 -516
<< ndiff >>
rect 206 -2621 264 -2609
rect 206 -2997 218 -2621
rect 252 -2997 264 -2621
rect 206 -3009 264 -2997
rect 294 -2621 352 -2609
rect 294 -2997 306 -2621
rect 340 -2997 352 -2621
rect 294 -3009 352 -2997
rect 486 -2621 544 -2609
rect 486 -2997 498 -2621
rect 532 -2997 544 -2621
rect 486 -3009 544 -2997
rect 574 -2621 632 -2609
rect 574 -2997 586 -2621
rect 620 -2997 632 -2621
rect 574 -3009 632 -2997
rect 766 -2621 824 -2609
rect 766 -2997 778 -2621
rect 812 -2997 824 -2621
rect 766 -3009 824 -2997
rect 854 -2621 912 -2609
rect 854 -2997 866 -2621
rect 900 -2997 912 -2621
rect 854 -3009 912 -2997
rect 1046 -2621 1104 -2609
rect 1046 -2997 1058 -2621
rect 1092 -2997 1104 -2621
rect 1046 -3009 1104 -2997
rect 1134 -2621 1192 -2609
rect 1134 -2997 1146 -2621
rect 1180 -2997 1192 -2621
rect 1134 -3009 1192 -2997
rect 1326 -2621 1384 -2609
rect 1326 -2997 1338 -2621
rect 1372 -2997 1384 -2621
rect 1326 -3009 1384 -2997
rect 1414 -2621 1472 -2609
rect 1414 -2997 1426 -2621
rect 1460 -2997 1472 -2621
rect 1414 -3009 1472 -2997
rect 1606 -2621 1664 -2609
rect 1606 -2997 1618 -2621
rect 1652 -2997 1664 -2621
rect 1606 -3009 1664 -2997
rect 1694 -2621 1752 -2609
rect 1694 -2997 1706 -2621
rect 1740 -2997 1752 -2621
rect 1694 -3009 1752 -2997
rect 1886 -2621 1944 -2609
rect 1886 -2997 1898 -2621
rect 1932 -2997 1944 -2621
rect 1886 -3009 1944 -2997
rect 1974 -2621 2032 -2609
rect 1974 -2997 1986 -2621
rect 2020 -2997 2032 -2621
rect 1974 -3009 2032 -2997
rect 2166 -2621 2224 -2609
rect 2166 -2997 2178 -2621
rect 2212 -2997 2224 -2621
rect 2166 -3009 2224 -2997
rect 2254 -2621 2312 -2609
rect 2254 -2997 2266 -2621
rect 2300 -2997 2312 -2621
rect 2254 -3009 2312 -2997
rect 2446 -2621 2504 -2609
rect 2446 -2997 2458 -2621
rect 2492 -2997 2504 -2621
rect 2446 -3009 2504 -2997
rect 2534 -2621 2592 -2609
rect 2534 -2997 2546 -2621
rect 2580 -2997 2592 -2621
rect 2534 -3009 2592 -2997
rect 2726 -2621 2784 -2609
rect 2726 -2997 2738 -2621
rect 2772 -2997 2784 -2621
rect 2726 -3009 2784 -2997
rect 2814 -2621 2872 -2609
rect 2814 -2997 2826 -2621
rect 2860 -2997 2872 -2621
rect 2814 -3009 2872 -2997
rect 206 -3441 264 -3429
rect 206 -3817 218 -3441
rect 252 -3817 264 -3441
rect 206 -3829 264 -3817
rect 294 -3441 352 -3429
rect 294 -3817 306 -3441
rect 340 -3817 352 -3441
rect 294 -3829 352 -3817
rect 486 -3441 544 -3429
rect 486 -3817 498 -3441
rect 532 -3817 544 -3441
rect 486 -3829 544 -3817
rect 574 -3441 632 -3429
rect 574 -3817 586 -3441
rect 620 -3817 632 -3441
rect 574 -3829 632 -3817
rect 766 -3441 824 -3429
rect 766 -3817 778 -3441
rect 812 -3817 824 -3441
rect 766 -3829 824 -3817
rect 854 -3441 912 -3429
rect 854 -3817 866 -3441
rect 900 -3817 912 -3441
rect 854 -3829 912 -3817
rect 1046 -3441 1104 -3429
rect 1046 -3817 1058 -3441
rect 1092 -3817 1104 -3441
rect 1046 -3829 1104 -3817
rect 1134 -3441 1192 -3429
rect 1134 -3817 1146 -3441
rect 1180 -3817 1192 -3441
rect 1134 -3829 1192 -3817
rect 1326 -3441 1384 -3429
rect 1326 -3817 1338 -3441
rect 1372 -3817 1384 -3441
rect 1326 -3829 1384 -3817
rect 1414 -3441 1472 -3429
rect 1414 -3817 1426 -3441
rect 1460 -3817 1472 -3441
rect 1414 -3829 1472 -3817
rect 1606 -3441 1664 -3429
rect 1606 -3817 1618 -3441
rect 1652 -3817 1664 -3441
rect 1606 -3829 1664 -3817
rect 1694 -3441 1752 -3429
rect 1694 -3817 1706 -3441
rect 1740 -3817 1752 -3441
rect 1694 -3829 1752 -3817
rect 1886 -3441 1944 -3429
rect 1886 -3817 1898 -3441
rect 1932 -3817 1944 -3441
rect 1886 -3829 1944 -3817
rect 1974 -3441 2032 -3429
rect 1974 -3817 1986 -3441
rect 2020 -3817 2032 -3441
rect 1974 -3829 2032 -3817
rect 2166 -3441 2224 -3429
rect 2166 -3817 2178 -3441
rect 2212 -3817 2224 -3441
rect 2166 -3829 2224 -3817
rect 2254 -3441 2312 -3429
rect 2254 -3817 2266 -3441
rect 2300 -3817 2312 -3441
rect 2254 -3829 2312 -3817
rect 2446 -3441 2504 -3429
rect 2446 -3817 2458 -3441
rect 2492 -3817 2504 -3441
rect 2446 -3829 2504 -3817
rect 2534 -3441 2592 -3429
rect 2534 -3817 2546 -3441
rect 2580 -3817 2592 -3441
rect 2534 -3829 2592 -3817
rect 2726 -3441 2784 -3429
rect 2726 -3817 2738 -3441
rect 2772 -3817 2784 -3441
rect 2726 -3829 2784 -3817
rect 2814 -3441 2872 -3429
rect 2814 -3817 2826 -3441
rect 2860 -3817 2872 -3441
rect 2814 -3829 2872 -3817
rect 1326 -4721 1384 -4709
rect 1326 -5097 1338 -4721
rect 1372 -5097 1384 -4721
rect 1326 -5109 1384 -5097
rect 1414 -4721 1472 -4709
rect 1414 -5097 1426 -4721
rect 1460 -5097 1472 -4721
rect 1414 -5109 1472 -5097
rect 1606 -4721 1664 -4709
rect 1606 -5097 1618 -4721
rect 1652 -5097 1664 -4721
rect 1606 -5109 1664 -5097
rect 1694 -4721 1752 -4709
rect 1694 -5097 1706 -4721
rect 1740 -5097 1752 -4721
rect 1694 -5109 1752 -5097
rect 1325 -5579 1383 -5567
rect 1325 -5955 1337 -5579
rect 1371 -5955 1383 -5579
rect 1325 -5967 1383 -5955
rect 1413 -5579 1471 -5567
rect 1413 -5955 1425 -5579
rect 1459 -5955 1471 -5579
rect 1413 -5967 1471 -5955
rect 1605 -5579 1663 -5567
rect 1605 -5955 1617 -5579
rect 1651 -5955 1663 -5579
rect 1605 -5967 1663 -5955
rect 1693 -5579 1751 -5567
rect 1693 -5955 1705 -5579
rect 1739 -5955 1751 -5579
rect 1693 -5967 1751 -5955
rect 206 -6524 264 -6512
rect 206 -6900 218 -6524
rect 252 -6900 264 -6524
rect 206 -6912 264 -6900
rect 294 -6524 352 -6512
rect 294 -6900 306 -6524
rect 340 -6900 352 -6524
rect 294 -6912 352 -6900
rect 486 -6524 544 -6512
rect 486 -6900 498 -6524
rect 532 -6900 544 -6524
rect 486 -6912 544 -6900
rect 574 -6524 632 -6512
rect 574 -6900 586 -6524
rect 620 -6900 632 -6524
rect 574 -6912 632 -6900
rect 766 -6524 824 -6512
rect 766 -6900 778 -6524
rect 812 -6900 824 -6524
rect 766 -6912 824 -6900
rect 854 -6524 912 -6512
rect 854 -6900 866 -6524
rect 900 -6900 912 -6524
rect 854 -6912 912 -6900
rect 1046 -6524 1104 -6512
rect 1046 -6900 1058 -6524
rect 1092 -6900 1104 -6524
rect 1046 -6912 1104 -6900
rect 1134 -6524 1192 -6512
rect 1134 -6900 1146 -6524
rect 1180 -6900 1192 -6524
rect 1134 -6912 1192 -6900
rect 1326 -6524 1384 -6512
rect 1326 -6900 1338 -6524
rect 1372 -6900 1384 -6524
rect 1326 -6912 1384 -6900
rect 1414 -6524 1472 -6512
rect 1414 -6900 1426 -6524
rect 1460 -6900 1472 -6524
rect 1414 -6912 1472 -6900
rect 1606 -6524 1664 -6512
rect 1606 -6900 1618 -6524
rect 1652 -6900 1664 -6524
rect 1606 -6912 1664 -6900
rect 1694 -6524 1752 -6512
rect 1694 -6900 1706 -6524
rect 1740 -6900 1752 -6524
rect 1694 -6912 1752 -6900
rect 1886 -6524 1944 -6512
rect 1886 -6900 1898 -6524
rect 1932 -6900 1944 -6524
rect 1886 -6912 1944 -6900
rect 1974 -6524 2032 -6512
rect 1974 -6900 1986 -6524
rect 2020 -6900 2032 -6524
rect 1974 -6912 2032 -6900
rect 2166 -6524 2224 -6512
rect 2166 -6900 2178 -6524
rect 2212 -6900 2224 -6524
rect 2166 -6912 2224 -6900
rect 2254 -6524 2312 -6512
rect 2254 -6900 2266 -6524
rect 2300 -6900 2312 -6524
rect 2254 -6912 2312 -6900
rect 2446 -6524 2504 -6512
rect 2446 -6900 2458 -6524
rect 2492 -6900 2504 -6524
rect 2446 -6912 2504 -6900
rect 2534 -6524 2592 -6512
rect 2534 -6900 2546 -6524
rect 2580 -6900 2592 -6524
rect 2534 -6912 2592 -6900
rect 2726 -6524 2784 -6512
rect 2726 -6900 2738 -6524
rect 2772 -6900 2784 -6524
rect 2726 -6912 2784 -6900
rect 2814 -6524 2872 -6512
rect 2814 -6900 2826 -6524
rect 2860 -6900 2872 -6524
rect 2814 -6912 2872 -6900
rect 206 -7222 264 -7210
rect 206 -7598 218 -7222
rect 252 -7598 264 -7222
rect 206 -7610 264 -7598
rect 294 -7222 352 -7210
rect 294 -7598 306 -7222
rect 340 -7598 352 -7222
rect 294 -7610 352 -7598
rect 486 -7222 544 -7210
rect 486 -7598 498 -7222
rect 532 -7598 544 -7222
rect 486 -7610 544 -7598
rect 574 -7222 632 -7210
rect 574 -7598 586 -7222
rect 620 -7598 632 -7222
rect 574 -7610 632 -7598
rect 766 -7222 824 -7210
rect 766 -7598 778 -7222
rect 812 -7598 824 -7222
rect 766 -7610 824 -7598
rect 854 -7222 912 -7210
rect 854 -7598 866 -7222
rect 900 -7598 912 -7222
rect 854 -7610 912 -7598
rect 1046 -7222 1104 -7210
rect 1046 -7598 1058 -7222
rect 1092 -7598 1104 -7222
rect 1046 -7610 1104 -7598
rect 1134 -7222 1192 -7210
rect 1134 -7598 1146 -7222
rect 1180 -7598 1192 -7222
rect 1134 -7610 1192 -7598
rect 1326 -7222 1384 -7210
rect 1326 -7598 1338 -7222
rect 1372 -7598 1384 -7222
rect 1326 -7610 1384 -7598
rect 1414 -7222 1472 -7210
rect 1414 -7598 1426 -7222
rect 1460 -7598 1472 -7222
rect 1414 -7610 1472 -7598
rect 1606 -7222 1664 -7210
rect 1606 -7598 1618 -7222
rect 1652 -7598 1664 -7222
rect 1606 -7610 1664 -7598
rect 1694 -7222 1752 -7210
rect 1694 -7598 1706 -7222
rect 1740 -7598 1752 -7222
rect 1694 -7610 1752 -7598
rect 1886 -7222 1944 -7210
rect 1886 -7598 1898 -7222
rect 1932 -7598 1944 -7222
rect 1886 -7610 1944 -7598
rect 1974 -7222 2032 -7210
rect 1974 -7598 1986 -7222
rect 2020 -7598 2032 -7222
rect 1974 -7610 2032 -7598
rect 2166 -7222 2224 -7210
rect 2166 -7598 2178 -7222
rect 2212 -7598 2224 -7222
rect 2166 -7610 2224 -7598
rect 2254 -7222 2312 -7210
rect 2254 -7598 2266 -7222
rect 2300 -7598 2312 -7222
rect 2254 -7610 2312 -7598
rect 2446 -7222 2504 -7210
rect 2446 -7598 2458 -7222
rect 2492 -7598 2504 -7222
rect 2446 -7610 2504 -7598
rect 2534 -7222 2592 -7210
rect 2534 -7598 2546 -7222
rect 2580 -7598 2592 -7222
rect 2534 -7610 2592 -7598
rect 2726 -7222 2784 -7210
rect 2726 -7598 2738 -7222
rect 2772 -7598 2784 -7222
rect 2726 -7610 2784 -7598
rect 2814 -7222 2872 -7210
rect 2814 -7598 2826 -7222
rect 2860 -7598 2872 -7222
rect 2814 -7610 2872 -7598
<< pdiff >>
rect -73 188 -15 200
rect -73 -188 -61 188
rect -27 -188 -15 188
rect -73 -200 -15 -188
rect 15 188 73 200
rect 15 -188 27 188
rect 61 -188 73 188
rect 15 -200 73 -188
rect 207 188 265 200
rect 207 -188 219 188
rect 253 -188 265 188
rect 207 -200 265 -188
rect 295 188 353 200
rect 295 -188 307 188
rect 341 -188 353 188
rect 295 -200 353 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 575 188 633 200
rect 575 -188 587 188
rect 621 -188 633 188
rect 575 -200 633 -188
rect 767 188 825 200
rect 767 -188 779 188
rect 813 -188 825 188
rect 767 -200 825 -188
rect 855 188 913 200
rect 855 -188 867 188
rect 901 -188 913 188
rect 855 -200 913 -188
rect 1047 188 1105 200
rect 1047 -188 1059 188
rect 1093 -188 1105 188
rect 1047 -200 1105 -188
rect 1135 188 1193 200
rect 1135 -188 1147 188
rect 1181 -188 1193 188
rect 1135 -200 1193 -188
rect 1327 188 1385 200
rect 1327 -188 1339 188
rect 1373 -188 1385 188
rect 1327 -200 1385 -188
rect 1415 188 1473 200
rect 1415 -188 1427 188
rect 1461 -188 1473 188
rect 1415 -200 1473 -188
rect 1607 188 1665 200
rect 1607 -188 1619 188
rect 1653 -188 1665 188
rect 1607 -200 1665 -188
rect 1695 188 1753 200
rect 1695 -188 1707 188
rect 1741 -188 1753 188
rect 1695 -200 1753 -188
rect 1887 188 1945 200
rect 1887 -188 1899 188
rect 1933 -188 1945 188
rect 1887 -200 1945 -188
rect 1975 188 2033 200
rect 1975 -188 1987 188
rect 2021 -188 2033 188
rect 1975 -200 2033 -188
rect 2167 188 2225 200
rect 2167 -188 2179 188
rect 2213 -188 2225 188
rect 2167 -200 2225 -188
rect 2255 188 2313 200
rect 2255 -188 2267 188
rect 2301 -188 2313 188
rect 2255 -200 2313 -188
rect 2447 188 2505 200
rect 2447 -188 2459 188
rect 2493 -188 2505 188
rect 2447 -200 2505 -188
rect 2535 188 2593 200
rect 2535 -188 2547 188
rect 2581 -188 2593 188
rect 2535 -200 2593 -188
rect 2727 188 2785 200
rect 2727 -188 2739 188
rect 2773 -188 2785 188
rect 2727 -200 2785 -188
rect 2815 188 2873 200
rect 2815 -188 2827 188
rect 2861 -188 2873 188
rect 2815 -200 2873 -188
rect 3007 188 3065 200
rect 3007 -188 3019 188
rect 3053 -188 3065 188
rect 3007 -200 3065 -188
rect 3095 188 3153 200
rect 3095 -188 3107 188
rect 3141 -188 3153 188
rect 3095 -200 3153 -188
rect -73 -528 -15 -516
rect -73 -904 -61 -528
rect -27 -904 -15 -528
rect -73 -916 -15 -904
rect 15 -528 73 -516
rect 15 -904 27 -528
rect 61 -904 73 -528
rect 15 -916 73 -904
rect 207 -528 265 -516
rect 207 -904 219 -528
rect 253 -904 265 -528
rect 207 -916 265 -904
rect 295 -528 353 -516
rect 295 -904 307 -528
rect 341 -904 353 -528
rect 295 -916 353 -904
rect 487 -528 545 -516
rect 487 -904 499 -528
rect 533 -904 545 -528
rect 487 -916 545 -904
rect 575 -528 633 -516
rect 575 -904 587 -528
rect 621 -904 633 -528
rect 575 -916 633 -904
rect 767 -528 825 -516
rect 767 -904 779 -528
rect 813 -904 825 -528
rect 767 -916 825 -904
rect 855 -528 913 -516
rect 855 -904 867 -528
rect 901 -904 913 -528
rect 855 -916 913 -904
rect 1047 -528 1105 -516
rect 1047 -904 1059 -528
rect 1093 -904 1105 -528
rect 1047 -916 1105 -904
rect 1135 -528 1193 -516
rect 1135 -904 1147 -528
rect 1181 -904 1193 -528
rect 1135 -916 1193 -904
rect 1327 -528 1385 -516
rect 1327 -904 1339 -528
rect 1373 -904 1385 -528
rect 1327 -916 1385 -904
rect 1415 -528 1473 -516
rect 1415 -904 1427 -528
rect 1461 -904 1473 -528
rect 1415 -916 1473 -904
rect 1607 -528 1665 -516
rect 1607 -904 1619 -528
rect 1653 -904 1665 -528
rect 1607 -916 1665 -904
rect 1695 -528 1753 -516
rect 1695 -904 1707 -528
rect 1741 -904 1753 -528
rect 1695 -916 1753 -904
rect 1887 -528 1945 -516
rect 1887 -904 1899 -528
rect 1933 -904 1945 -528
rect 1887 -916 1945 -904
rect 1975 -528 2033 -516
rect 1975 -904 1987 -528
rect 2021 -904 2033 -528
rect 1975 -916 2033 -904
rect 2167 -528 2225 -516
rect 2167 -904 2179 -528
rect 2213 -904 2225 -528
rect 2167 -916 2225 -904
rect 2255 -528 2313 -516
rect 2255 -904 2267 -528
rect 2301 -904 2313 -528
rect 2255 -916 2313 -904
rect 2447 -528 2505 -516
rect 2447 -904 2459 -528
rect 2493 -904 2505 -528
rect 2447 -916 2505 -904
rect 2535 -528 2593 -516
rect 2535 -904 2547 -528
rect 2581 -904 2593 -528
rect 2535 -916 2593 -904
rect 2727 -528 2785 -516
rect 2727 -904 2739 -528
rect 2773 -904 2785 -528
rect 2727 -916 2785 -904
rect 2815 -528 2873 -516
rect 2815 -904 2827 -528
rect 2861 -904 2873 -528
rect 2815 -916 2873 -904
rect 3007 -528 3065 -516
rect 3007 -904 3019 -528
rect 3053 -904 3065 -528
rect 3007 -916 3065 -904
rect 3095 -528 3153 -516
rect 3095 -904 3107 -528
rect 3141 -904 3153 -528
rect 3095 -916 3153 -904
<< ndiffc >>
rect 218 -2997 252 -2621
rect 306 -2997 340 -2621
rect 498 -2997 532 -2621
rect 586 -2997 620 -2621
rect 778 -2997 812 -2621
rect 866 -2997 900 -2621
rect 1058 -2997 1092 -2621
rect 1146 -2997 1180 -2621
rect 1338 -2997 1372 -2621
rect 1426 -2997 1460 -2621
rect 1618 -2997 1652 -2621
rect 1706 -2997 1740 -2621
rect 1898 -2997 1932 -2621
rect 1986 -2997 2020 -2621
rect 2178 -2997 2212 -2621
rect 2266 -2997 2300 -2621
rect 2458 -2997 2492 -2621
rect 2546 -2997 2580 -2621
rect 2738 -2997 2772 -2621
rect 2826 -2997 2860 -2621
rect 218 -3817 252 -3441
rect 306 -3817 340 -3441
rect 498 -3817 532 -3441
rect 586 -3817 620 -3441
rect 778 -3817 812 -3441
rect 866 -3817 900 -3441
rect 1058 -3817 1092 -3441
rect 1146 -3817 1180 -3441
rect 1338 -3817 1372 -3441
rect 1426 -3817 1460 -3441
rect 1618 -3817 1652 -3441
rect 1706 -3817 1740 -3441
rect 1898 -3817 1932 -3441
rect 1986 -3817 2020 -3441
rect 2178 -3817 2212 -3441
rect 2266 -3817 2300 -3441
rect 2458 -3817 2492 -3441
rect 2546 -3817 2580 -3441
rect 2738 -3817 2772 -3441
rect 2826 -3817 2860 -3441
rect 1338 -5097 1372 -4721
rect 1426 -5097 1460 -4721
rect 1618 -5097 1652 -4721
rect 1706 -5097 1740 -4721
rect 1337 -5955 1371 -5579
rect 1425 -5955 1459 -5579
rect 1617 -5955 1651 -5579
rect 1705 -5955 1739 -5579
rect 218 -6900 252 -6524
rect 306 -6900 340 -6524
rect 498 -6900 532 -6524
rect 586 -6900 620 -6524
rect 778 -6900 812 -6524
rect 866 -6900 900 -6524
rect 1058 -6900 1092 -6524
rect 1146 -6900 1180 -6524
rect 1338 -6900 1372 -6524
rect 1426 -6900 1460 -6524
rect 1618 -6900 1652 -6524
rect 1706 -6900 1740 -6524
rect 1898 -6900 1932 -6524
rect 1986 -6900 2020 -6524
rect 2178 -6900 2212 -6524
rect 2266 -6900 2300 -6524
rect 2458 -6900 2492 -6524
rect 2546 -6900 2580 -6524
rect 2738 -6900 2772 -6524
rect 2826 -6900 2860 -6524
rect 218 -7598 252 -7222
rect 306 -7598 340 -7222
rect 498 -7598 532 -7222
rect 586 -7598 620 -7222
rect 778 -7598 812 -7222
rect 866 -7598 900 -7222
rect 1058 -7598 1092 -7222
rect 1146 -7598 1180 -7222
rect 1338 -7598 1372 -7222
rect 1426 -7598 1460 -7222
rect 1618 -7598 1652 -7222
rect 1706 -7598 1740 -7222
rect 1898 -7598 1932 -7222
rect 1986 -7598 2020 -7222
rect 2178 -7598 2212 -7222
rect 2266 -7598 2300 -7222
rect 2458 -7598 2492 -7222
rect 2546 -7598 2580 -7222
rect 2738 -7598 2772 -7222
rect 2826 -7598 2860 -7222
<< pdiffc >>
rect -61 -188 -27 188
rect 27 -188 61 188
rect 219 -188 253 188
rect 307 -188 341 188
rect 499 -188 533 188
rect 587 -188 621 188
rect 779 -188 813 188
rect 867 -188 901 188
rect 1059 -188 1093 188
rect 1147 -188 1181 188
rect 1339 -188 1373 188
rect 1427 -188 1461 188
rect 1619 -188 1653 188
rect 1707 -188 1741 188
rect 1899 -188 1933 188
rect 1987 -188 2021 188
rect 2179 -188 2213 188
rect 2267 -188 2301 188
rect 2459 -188 2493 188
rect 2547 -188 2581 188
rect 2739 -188 2773 188
rect 2827 -188 2861 188
rect 3019 -188 3053 188
rect 3107 -188 3141 188
rect -61 -904 -27 -528
rect 27 -904 61 -528
rect 219 -904 253 -528
rect 307 -904 341 -528
rect 499 -904 533 -528
rect 587 -904 621 -528
rect 779 -904 813 -528
rect 867 -904 901 -528
rect 1059 -904 1093 -528
rect 1147 -904 1181 -528
rect 1339 -904 1373 -528
rect 1427 -904 1461 -528
rect 1619 -904 1653 -528
rect 1707 -904 1741 -528
rect 1899 -904 1933 -528
rect 1987 -904 2021 -528
rect 2179 -904 2213 -528
rect 2267 -904 2301 -528
rect 2459 -904 2493 -528
rect 2547 -904 2581 -528
rect 2739 -904 2773 -528
rect 2827 -904 2861 -528
rect 3019 -904 3053 -528
rect 3107 -904 3141 -528
<< mvpsubdiff >>
rect -508 -1978 3746 -1966
rect -508 -2078 -334 -1978
rect 3572 -2078 3746 -1978
rect -508 -2090 3746 -2078
rect -508 -2140 -384 -2090
rect -508 -8432 -496 -2140
rect -396 -8432 -384 -2140
rect 3622 -2140 3746 -2090
rect -508 -8482 -384 -8432
rect 3622 -8432 3634 -2140
rect 3734 -8432 3746 -2140
rect 3622 -8482 3746 -8432
rect -508 -8494 3746 -8482
rect -508 -8594 -334 -8494
rect 3572 -8594 3746 -8494
rect -508 -8606 3746 -8594
<< mvnsubdiff >>
rect -508 1122 3746 1134
rect -508 1022 -334 1122
rect 3572 1022 3746 1122
rect -508 1010 3746 1022
rect -508 960 -384 1010
rect -508 -1540 -496 960
rect -396 -1540 -384 960
rect 3622 960 3746 1010
rect -508 -1590 -384 -1540
rect 3622 -1540 3634 960
rect 3734 -1540 3746 960
rect 3622 -1590 3746 -1540
rect -508 -1602 3746 -1590
rect -508 -1702 -334 -1602
rect 3572 -1702 3746 -1602
rect -508 -1714 3746 -1702
<< mvpsubdiffcont >>
rect -334 -2078 3572 -1978
rect -496 -8432 -396 -2140
rect 3634 -8432 3734 -2140
rect -334 -8594 3572 -8494
<< mvnsubdiffcont >>
rect -334 1022 3572 1122
rect -496 -1540 -396 960
rect 3634 -1540 3734 960
rect -334 -1702 3572 -1602
<< poly >>
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect 247 281 313 297
rect 247 247 263 281
rect 297 247 313 281
rect 247 231 313 247
rect 527 281 593 297
rect 527 247 543 281
rect 577 247 593 281
rect 527 231 593 247
rect 807 281 873 297
rect 807 247 823 281
rect 857 247 873 281
rect 807 231 873 247
rect 1087 281 1153 297
rect 1087 247 1103 281
rect 1137 247 1153 281
rect 1087 231 1153 247
rect 1367 281 1433 297
rect 1367 247 1383 281
rect 1417 247 1433 281
rect 1367 231 1433 247
rect 1647 281 1713 297
rect 1647 247 1663 281
rect 1697 247 1713 281
rect 1647 231 1713 247
rect 1927 281 1993 297
rect 1927 247 1943 281
rect 1977 247 1993 281
rect 1927 231 1993 247
rect 2207 281 2273 297
rect 2207 247 2223 281
rect 2257 247 2273 281
rect 2207 231 2273 247
rect 2487 281 2553 297
rect 2487 247 2503 281
rect 2537 247 2553 281
rect 2487 231 2553 247
rect 2767 281 2833 297
rect 2767 247 2783 281
rect 2817 247 2833 281
rect 2767 231 2833 247
rect 3047 281 3113 297
rect 3047 247 3063 281
rect 3097 247 3113 281
rect 3047 231 3113 247
rect -15 200 15 231
rect 265 200 295 231
rect 545 200 575 231
rect 825 200 855 231
rect 1105 200 1135 231
rect 1385 200 1415 231
rect 1665 200 1695 231
rect 1945 200 1975 231
rect 2225 200 2255 231
rect 2505 200 2535 231
rect 2785 200 2815 231
rect 3065 200 3095 231
rect -15 -231 15 -200
rect 265 -231 295 -200
rect 545 -231 575 -200
rect 825 -231 855 -200
rect 1105 -231 1135 -200
rect 1385 -231 1415 -200
rect 1665 -231 1695 -200
rect 1945 -231 1975 -200
rect 2225 -231 2255 -200
rect 2505 -231 2535 -200
rect 2785 -231 2815 -200
rect 3065 -231 3095 -200
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
rect 247 -247 313 -231
rect 247 -281 263 -247
rect 297 -281 313 -247
rect 247 -297 313 -281
rect 527 -247 593 -231
rect 527 -281 543 -247
rect 577 -281 593 -247
rect 527 -297 593 -281
rect 807 -247 873 -231
rect 807 -281 823 -247
rect 857 -281 873 -247
rect 807 -297 873 -281
rect 1087 -247 1153 -231
rect 1087 -281 1103 -247
rect 1137 -281 1153 -247
rect 1087 -297 1153 -281
rect 1367 -247 1433 -231
rect 1367 -281 1383 -247
rect 1417 -281 1433 -247
rect 1367 -297 1433 -281
rect 1647 -247 1713 -231
rect 1647 -281 1663 -247
rect 1697 -281 1713 -247
rect 1647 -297 1713 -281
rect 1927 -247 1993 -231
rect 1927 -281 1943 -247
rect 1977 -281 1993 -247
rect 1927 -297 1993 -281
rect 2207 -247 2273 -231
rect 2207 -281 2223 -247
rect 2257 -281 2273 -247
rect 2207 -297 2273 -281
rect 2487 -247 2553 -231
rect 2487 -281 2503 -247
rect 2537 -281 2553 -247
rect 2487 -297 2553 -281
rect 2767 -247 2833 -231
rect 2767 -281 2783 -247
rect 2817 -281 2833 -247
rect 2767 -297 2833 -281
rect 3047 -247 3113 -231
rect 3047 -281 3063 -247
rect 3097 -281 3113 -247
rect 3047 -297 3113 -281
rect -33 -435 33 -419
rect -33 -469 -17 -435
rect 17 -469 33 -435
rect -33 -485 33 -469
rect 247 -435 313 -419
rect 247 -469 263 -435
rect 297 -469 313 -435
rect 247 -485 313 -469
rect 527 -435 593 -419
rect 527 -469 543 -435
rect 577 -469 593 -435
rect 527 -485 593 -469
rect 807 -435 873 -419
rect 807 -469 823 -435
rect 857 -469 873 -435
rect 807 -485 873 -469
rect 1087 -435 1153 -419
rect 1087 -469 1103 -435
rect 1137 -469 1153 -435
rect 1087 -485 1153 -469
rect 1367 -435 1433 -419
rect 1367 -469 1383 -435
rect 1417 -469 1433 -435
rect 1367 -485 1433 -469
rect 1647 -435 1713 -419
rect 1647 -469 1663 -435
rect 1697 -469 1713 -435
rect 1647 -485 1713 -469
rect 1927 -435 1993 -419
rect 1927 -469 1943 -435
rect 1977 -469 1993 -435
rect 1927 -485 1993 -469
rect 2207 -435 2273 -419
rect 2207 -469 2223 -435
rect 2257 -469 2273 -435
rect 2207 -485 2273 -469
rect 2487 -435 2553 -419
rect 2487 -469 2503 -435
rect 2537 -469 2553 -435
rect 2487 -485 2553 -469
rect 2767 -435 2833 -419
rect 2767 -469 2783 -435
rect 2817 -469 2833 -435
rect 2767 -485 2833 -469
rect 3047 -435 3113 -419
rect 3047 -469 3063 -435
rect 3097 -469 3113 -435
rect 3047 -485 3113 -469
rect -15 -516 15 -485
rect 265 -516 295 -485
rect 545 -516 575 -485
rect 825 -516 855 -485
rect 1105 -516 1135 -485
rect 1385 -516 1415 -485
rect 1665 -516 1695 -485
rect 1945 -516 1975 -485
rect 2225 -516 2255 -485
rect 2505 -516 2535 -485
rect 2785 -516 2815 -485
rect 3065 -516 3095 -485
rect -15 -947 15 -916
rect 265 -947 295 -916
rect 545 -947 575 -916
rect 825 -947 855 -916
rect 1105 -947 1135 -916
rect 1385 -947 1415 -916
rect 1665 -947 1695 -916
rect 1945 -947 1975 -916
rect 2225 -947 2255 -916
rect 2505 -947 2535 -916
rect 2785 -947 2815 -916
rect 3065 -947 3095 -916
rect -33 -963 33 -947
rect -33 -997 -17 -963
rect 17 -997 33 -963
rect -33 -1013 33 -997
rect 247 -963 313 -947
rect 247 -997 263 -963
rect 297 -997 313 -963
rect 247 -1013 313 -997
rect 527 -963 593 -947
rect 527 -997 543 -963
rect 577 -997 593 -963
rect 527 -1013 593 -997
rect 807 -963 873 -947
rect 807 -997 823 -963
rect 857 -997 873 -963
rect 807 -1013 873 -997
rect 1087 -963 1153 -947
rect 1087 -997 1103 -963
rect 1137 -997 1153 -963
rect 1087 -1013 1153 -997
rect 1367 -963 1433 -947
rect 1367 -997 1383 -963
rect 1417 -997 1433 -963
rect 1367 -1013 1433 -997
rect 1647 -963 1713 -947
rect 1647 -997 1663 -963
rect 1697 -997 1713 -963
rect 1647 -1013 1713 -997
rect 1927 -963 1993 -947
rect 1927 -997 1943 -963
rect 1977 -997 1993 -963
rect 1927 -1013 1993 -997
rect 2207 -963 2273 -947
rect 2207 -997 2223 -963
rect 2257 -997 2273 -963
rect 2207 -1013 2273 -997
rect 2487 -963 2553 -947
rect 2487 -997 2503 -963
rect 2537 -997 2553 -963
rect 2487 -1013 2553 -997
rect 2767 -963 2833 -947
rect 2767 -997 2783 -963
rect 2817 -997 2833 -963
rect 2767 -1013 2833 -997
rect 3047 -963 3113 -947
rect 3047 -997 3063 -963
rect 3097 -997 3113 -963
rect 3047 -1013 3113 -997
rect 246 -2537 312 -2521
rect 246 -2571 262 -2537
rect 296 -2571 312 -2537
rect 246 -2587 312 -2571
rect 526 -2537 592 -2521
rect 526 -2571 542 -2537
rect 576 -2571 592 -2537
rect 526 -2587 592 -2571
rect 806 -2537 872 -2521
rect 806 -2571 822 -2537
rect 856 -2571 872 -2537
rect 806 -2587 872 -2571
rect 1086 -2537 1152 -2521
rect 1086 -2571 1102 -2537
rect 1136 -2571 1152 -2537
rect 1086 -2587 1152 -2571
rect 1366 -2537 1432 -2521
rect 1366 -2571 1382 -2537
rect 1416 -2571 1432 -2537
rect 1366 -2587 1432 -2571
rect 1646 -2537 1712 -2521
rect 1646 -2571 1662 -2537
rect 1696 -2571 1712 -2537
rect 1646 -2587 1712 -2571
rect 1926 -2537 1992 -2521
rect 1926 -2571 1942 -2537
rect 1976 -2571 1992 -2537
rect 1926 -2587 1992 -2571
rect 2206 -2537 2272 -2521
rect 2206 -2571 2222 -2537
rect 2256 -2571 2272 -2537
rect 2206 -2587 2272 -2571
rect 2486 -2537 2552 -2521
rect 2486 -2571 2502 -2537
rect 2536 -2571 2552 -2537
rect 2486 -2587 2552 -2571
rect 2766 -2537 2832 -2521
rect 2766 -2571 2782 -2537
rect 2816 -2571 2832 -2537
rect 2766 -2587 2832 -2571
rect 264 -2609 294 -2587
rect 544 -2609 574 -2587
rect 824 -2609 854 -2587
rect 1104 -2609 1134 -2587
rect 1384 -2609 1414 -2587
rect 1664 -2609 1694 -2587
rect 1944 -2609 1974 -2587
rect 2224 -2609 2254 -2587
rect 2504 -2609 2534 -2587
rect 2784 -2609 2814 -2587
rect 264 -3031 294 -3009
rect 544 -3031 574 -3009
rect 824 -3031 854 -3009
rect 1104 -3031 1134 -3009
rect 1384 -3031 1414 -3009
rect 1664 -3031 1694 -3009
rect 1944 -3031 1974 -3009
rect 2224 -3031 2254 -3009
rect 2504 -3031 2534 -3009
rect 2784 -3031 2814 -3009
rect 246 -3047 312 -3031
rect 246 -3081 262 -3047
rect 296 -3081 312 -3047
rect 246 -3097 312 -3081
rect 526 -3047 592 -3031
rect 526 -3081 542 -3047
rect 576 -3081 592 -3047
rect 526 -3097 592 -3081
rect 806 -3047 872 -3031
rect 806 -3081 822 -3047
rect 856 -3081 872 -3047
rect 806 -3097 872 -3081
rect 1086 -3047 1152 -3031
rect 1086 -3081 1102 -3047
rect 1136 -3081 1152 -3047
rect 1086 -3097 1152 -3081
rect 1366 -3047 1432 -3031
rect 1366 -3081 1382 -3047
rect 1416 -3081 1432 -3047
rect 1366 -3097 1432 -3081
rect 1646 -3047 1712 -3031
rect 1646 -3081 1662 -3047
rect 1696 -3081 1712 -3047
rect 1646 -3097 1712 -3081
rect 1926 -3047 1992 -3031
rect 1926 -3081 1942 -3047
rect 1976 -3081 1992 -3047
rect 1926 -3097 1992 -3081
rect 2206 -3047 2272 -3031
rect 2206 -3081 2222 -3047
rect 2256 -3081 2272 -3047
rect 2206 -3097 2272 -3081
rect 2486 -3047 2552 -3031
rect 2486 -3081 2502 -3047
rect 2536 -3081 2552 -3047
rect 2486 -3097 2552 -3081
rect 2766 -3047 2832 -3031
rect 2766 -3081 2782 -3047
rect 2816 -3081 2832 -3047
rect 2766 -3097 2832 -3081
rect 246 -3357 312 -3341
rect 246 -3391 262 -3357
rect 296 -3391 312 -3357
rect 246 -3407 312 -3391
rect 526 -3357 592 -3341
rect 526 -3391 542 -3357
rect 576 -3391 592 -3357
rect 526 -3407 592 -3391
rect 806 -3357 872 -3341
rect 806 -3391 822 -3357
rect 856 -3391 872 -3357
rect 806 -3407 872 -3391
rect 1086 -3357 1152 -3341
rect 1086 -3391 1102 -3357
rect 1136 -3391 1152 -3357
rect 1086 -3407 1152 -3391
rect 1366 -3357 1432 -3341
rect 1366 -3391 1382 -3357
rect 1416 -3391 1432 -3357
rect 1366 -3407 1432 -3391
rect 1646 -3357 1712 -3341
rect 1646 -3391 1662 -3357
rect 1696 -3391 1712 -3357
rect 1646 -3407 1712 -3391
rect 1926 -3357 1992 -3341
rect 1926 -3391 1942 -3357
rect 1976 -3391 1992 -3357
rect 1926 -3407 1992 -3391
rect 2206 -3357 2272 -3341
rect 2206 -3391 2222 -3357
rect 2256 -3391 2272 -3357
rect 2206 -3407 2272 -3391
rect 2486 -3357 2552 -3341
rect 2486 -3391 2502 -3357
rect 2536 -3391 2552 -3357
rect 2486 -3407 2552 -3391
rect 2766 -3357 2832 -3341
rect 2766 -3391 2782 -3357
rect 2816 -3391 2832 -3357
rect 2766 -3407 2832 -3391
rect 264 -3429 294 -3407
rect 544 -3429 574 -3407
rect 824 -3429 854 -3407
rect 1104 -3429 1134 -3407
rect 1384 -3429 1414 -3407
rect 1664 -3429 1694 -3407
rect 1944 -3429 1974 -3407
rect 2224 -3429 2254 -3407
rect 2504 -3429 2534 -3407
rect 2784 -3429 2814 -3407
rect 264 -3851 294 -3829
rect 544 -3851 574 -3829
rect 824 -3851 854 -3829
rect 1104 -3851 1134 -3829
rect 1384 -3851 1414 -3829
rect 1664 -3851 1694 -3829
rect 1944 -3851 1974 -3829
rect 2224 -3851 2254 -3829
rect 2504 -3851 2534 -3829
rect 2784 -3851 2814 -3829
rect 246 -3867 312 -3851
rect 246 -3901 262 -3867
rect 296 -3901 312 -3867
rect 246 -3917 312 -3901
rect 526 -3867 592 -3851
rect 526 -3901 542 -3867
rect 576 -3901 592 -3867
rect 526 -3917 592 -3901
rect 806 -3867 872 -3851
rect 806 -3901 822 -3867
rect 856 -3901 872 -3867
rect 806 -3917 872 -3901
rect 1086 -3867 1152 -3851
rect 1086 -3901 1102 -3867
rect 1136 -3901 1152 -3867
rect 1086 -3917 1152 -3901
rect 1366 -3867 1432 -3851
rect 1366 -3901 1382 -3867
rect 1416 -3901 1432 -3867
rect 1366 -3917 1432 -3901
rect 1646 -3867 1712 -3851
rect 1646 -3901 1662 -3867
rect 1696 -3901 1712 -3867
rect 1646 -3917 1712 -3901
rect 1926 -3867 1992 -3851
rect 1926 -3901 1942 -3867
rect 1976 -3901 1992 -3867
rect 1926 -3917 1992 -3901
rect 2206 -3867 2272 -3851
rect 2206 -3901 2222 -3867
rect 2256 -3901 2272 -3867
rect 2206 -3917 2272 -3901
rect 2486 -3867 2552 -3851
rect 2486 -3901 2502 -3867
rect 2536 -3901 2552 -3867
rect 2486 -3917 2552 -3901
rect 2766 -3867 2832 -3851
rect 2766 -3901 2782 -3867
rect 2816 -3901 2832 -3867
rect 2766 -3917 2832 -3901
rect 1366 -4637 1432 -4621
rect 1366 -4671 1382 -4637
rect 1416 -4671 1432 -4637
rect 1366 -4687 1432 -4671
rect 1646 -4637 1712 -4621
rect 1646 -4671 1662 -4637
rect 1696 -4671 1712 -4637
rect 1646 -4687 1712 -4671
rect 1384 -4709 1414 -4687
rect 1664 -4709 1694 -4687
rect 1384 -5131 1414 -5109
rect 1664 -5131 1694 -5109
rect 1366 -5147 1432 -5131
rect 1366 -5181 1382 -5147
rect 1416 -5181 1432 -5147
rect 1366 -5197 1432 -5181
rect 1646 -5147 1712 -5131
rect 1646 -5181 1662 -5147
rect 1696 -5181 1712 -5147
rect 1646 -5197 1712 -5181
rect 1365 -5495 1431 -5479
rect 1365 -5529 1381 -5495
rect 1415 -5529 1431 -5495
rect 1365 -5545 1431 -5529
rect 1645 -5495 1711 -5479
rect 1645 -5529 1661 -5495
rect 1695 -5529 1711 -5495
rect 1645 -5545 1711 -5529
rect 1383 -5567 1413 -5545
rect 1663 -5567 1693 -5545
rect 1383 -5993 1413 -5967
rect 1663 -5993 1693 -5967
rect 246 -6440 312 -6424
rect 246 -6474 262 -6440
rect 296 -6474 312 -6440
rect 246 -6490 312 -6474
rect 526 -6440 592 -6424
rect 526 -6474 542 -6440
rect 576 -6474 592 -6440
rect 526 -6490 592 -6474
rect 806 -6440 872 -6424
rect 806 -6474 822 -6440
rect 856 -6474 872 -6440
rect 806 -6490 872 -6474
rect 1086 -6440 1152 -6424
rect 1086 -6474 1102 -6440
rect 1136 -6474 1152 -6440
rect 1086 -6490 1152 -6474
rect 1366 -6440 1432 -6424
rect 1366 -6474 1382 -6440
rect 1416 -6474 1432 -6440
rect 1366 -6490 1432 -6474
rect 1646 -6440 1712 -6424
rect 1646 -6474 1662 -6440
rect 1696 -6474 1712 -6440
rect 1646 -6490 1712 -6474
rect 1926 -6440 1992 -6424
rect 1926 -6474 1942 -6440
rect 1976 -6474 1992 -6440
rect 1926 -6490 1992 -6474
rect 2206 -6440 2272 -6424
rect 2206 -6474 2222 -6440
rect 2256 -6474 2272 -6440
rect 2206 -6490 2272 -6474
rect 2486 -6440 2552 -6424
rect 2486 -6474 2502 -6440
rect 2536 -6474 2552 -6440
rect 2486 -6490 2552 -6474
rect 2766 -6440 2832 -6424
rect 2766 -6474 2782 -6440
rect 2816 -6474 2832 -6440
rect 2766 -6490 2832 -6474
rect 264 -6512 294 -6490
rect 544 -6512 574 -6490
rect 824 -6512 854 -6490
rect 1104 -6512 1134 -6490
rect 1384 -6512 1414 -6490
rect 1664 -6512 1694 -6490
rect 1944 -6512 1974 -6490
rect 2224 -6512 2254 -6490
rect 2504 -6512 2534 -6490
rect 2784 -6512 2814 -6490
rect 264 -6938 294 -6912
rect 544 -6938 574 -6912
rect 824 -6938 854 -6912
rect 1104 -6938 1134 -6912
rect 1384 -6938 1414 -6912
rect 1664 -6938 1694 -6912
rect 1944 -6938 1974 -6912
rect 2224 -6938 2254 -6912
rect 2504 -6938 2534 -6912
rect 2784 -6938 2814 -6912
rect 264 -7210 294 -7184
rect 544 -7210 574 -7184
rect 824 -7210 854 -7184
rect 1104 -7210 1134 -7184
rect 1384 -7210 1414 -7184
rect 1664 -7210 1694 -7184
rect 1944 -7210 1974 -7184
rect 2224 -7210 2254 -7184
rect 2504 -7210 2534 -7184
rect 2784 -7210 2814 -7184
rect 264 -7632 294 -7610
rect 544 -7632 574 -7610
rect 824 -7632 854 -7610
rect 1104 -7632 1134 -7610
rect 1384 -7632 1414 -7610
rect 1664 -7632 1694 -7610
rect 1944 -7632 1974 -7610
rect 2224 -7632 2254 -7610
rect 2504 -7632 2534 -7610
rect 2784 -7632 2814 -7610
rect 246 -7648 312 -7632
rect 246 -7682 262 -7648
rect 296 -7682 312 -7648
rect 246 -7698 312 -7682
rect 526 -7648 592 -7632
rect 526 -7682 542 -7648
rect 576 -7682 592 -7648
rect 526 -7698 592 -7682
rect 806 -7648 872 -7632
rect 806 -7682 822 -7648
rect 856 -7682 872 -7648
rect 806 -7698 872 -7682
rect 1086 -7648 1152 -7632
rect 1086 -7682 1102 -7648
rect 1136 -7682 1152 -7648
rect 1086 -7698 1152 -7682
rect 1366 -7648 1432 -7632
rect 1366 -7682 1382 -7648
rect 1416 -7682 1432 -7648
rect 1366 -7698 1432 -7682
rect 1646 -7648 1712 -7632
rect 1646 -7682 1662 -7648
rect 1696 -7682 1712 -7648
rect 1646 -7698 1712 -7682
rect 1926 -7648 1992 -7632
rect 1926 -7682 1942 -7648
rect 1976 -7682 1992 -7648
rect 1926 -7698 1992 -7682
rect 2206 -7648 2272 -7632
rect 2206 -7682 2222 -7648
rect 2256 -7682 2272 -7648
rect 2206 -7698 2272 -7682
rect 2486 -7648 2552 -7632
rect 2486 -7682 2502 -7648
rect 2536 -7682 2552 -7648
rect 2486 -7698 2552 -7682
rect 2766 -7648 2832 -7632
rect 2766 -7682 2782 -7648
rect 2816 -7682 2832 -7648
rect 2766 -7698 2832 -7682
<< polycont >>
rect -17 247 17 281
rect 263 247 297 281
rect 543 247 577 281
rect 823 247 857 281
rect 1103 247 1137 281
rect 1383 247 1417 281
rect 1663 247 1697 281
rect 1943 247 1977 281
rect 2223 247 2257 281
rect 2503 247 2537 281
rect 2783 247 2817 281
rect 3063 247 3097 281
rect -17 -281 17 -247
rect 263 -281 297 -247
rect 543 -281 577 -247
rect 823 -281 857 -247
rect 1103 -281 1137 -247
rect 1383 -281 1417 -247
rect 1663 -281 1697 -247
rect 1943 -281 1977 -247
rect 2223 -281 2257 -247
rect 2503 -281 2537 -247
rect 2783 -281 2817 -247
rect 3063 -281 3097 -247
rect -17 -469 17 -435
rect 263 -469 297 -435
rect 543 -469 577 -435
rect 823 -469 857 -435
rect 1103 -469 1137 -435
rect 1383 -469 1417 -435
rect 1663 -469 1697 -435
rect 1943 -469 1977 -435
rect 2223 -469 2257 -435
rect 2503 -469 2537 -435
rect 2783 -469 2817 -435
rect 3063 -469 3097 -435
rect -17 -997 17 -963
rect 263 -997 297 -963
rect 543 -997 577 -963
rect 823 -997 857 -963
rect 1103 -997 1137 -963
rect 1383 -997 1417 -963
rect 1663 -997 1697 -963
rect 1943 -997 1977 -963
rect 2223 -997 2257 -963
rect 2503 -997 2537 -963
rect 2783 -997 2817 -963
rect 3063 -997 3097 -963
rect 262 -2571 296 -2537
rect 542 -2571 576 -2537
rect 822 -2571 856 -2537
rect 1102 -2571 1136 -2537
rect 1382 -2571 1416 -2537
rect 1662 -2571 1696 -2537
rect 1942 -2571 1976 -2537
rect 2222 -2571 2256 -2537
rect 2502 -2571 2536 -2537
rect 2782 -2571 2816 -2537
rect 262 -3081 296 -3047
rect 542 -3081 576 -3047
rect 822 -3081 856 -3047
rect 1102 -3081 1136 -3047
rect 1382 -3081 1416 -3047
rect 1662 -3081 1696 -3047
rect 1942 -3081 1976 -3047
rect 2222 -3081 2256 -3047
rect 2502 -3081 2536 -3047
rect 2782 -3081 2816 -3047
rect 262 -3391 296 -3357
rect 542 -3391 576 -3357
rect 822 -3391 856 -3357
rect 1102 -3391 1136 -3357
rect 1382 -3391 1416 -3357
rect 1662 -3391 1696 -3357
rect 1942 -3391 1976 -3357
rect 2222 -3391 2256 -3357
rect 2502 -3391 2536 -3357
rect 2782 -3391 2816 -3357
rect 262 -3901 296 -3867
rect 542 -3901 576 -3867
rect 822 -3901 856 -3867
rect 1102 -3901 1136 -3867
rect 1382 -3901 1416 -3867
rect 1662 -3901 1696 -3867
rect 1942 -3901 1976 -3867
rect 2222 -3901 2256 -3867
rect 2502 -3901 2536 -3867
rect 2782 -3901 2816 -3867
rect 1382 -4671 1416 -4637
rect 1662 -4671 1696 -4637
rect 1382 -5181 1416 -5147
rect 1662 -5181 1696 -5147
rect 1381 -5529 1415 -5495
rect 1661 -5529 1695 -5495
rect 262 -6474 296 -6440
rect 542 -6474 576 -6440
rect 822 -6474 856 -6440
rect 1102 -6474 1136 -6440
rect 1382 -6474 1416 -6440
rect 1662 -6474 1696 -6440
rect 1942 -6474 1976 -6440
rect 2222 -6474 2256 -6440
rect 2502 -6474 2536 -6440
rect 2782 -6474 2816 -6440
rect 262 -7682 296 -7648
rect 542 -7682 576 -7648
rect 822 -7682 856 -7648
rect 1102 -7682 1136 -7648
rect 1382 -7682 1416 -7648
rect 1662 -7682 1696 -7648
rect 1942 -7682 1976 -7648
rect 2222 -7682 2256 -7648
rect 2502 -7682 2536 -7648
rect 2782 -7682 2816 -7648
<< locali >>
rect -496 960 -396 1122
rect 3634 960 3734 1122
rect -33 247 -17 281
rect 17 247 33 281
rect 247 247 263 281
rect 297 247 313 281
rect 527 247 543 281
rect 577 247 593 281
rect 807 247 823 281
rect 857 247 873 281
rect 1087 247 1103 281
rect 1137 247 1153 281
rect 1367 247 1383 281
rect 1417 247 1433 281
rect 1647 247 1663 281
rect 1697 247 1713 281
rect 1927 247 1943 281
rect 1977 247 1993 281
rect 2207 247 2223 281
rect 2257 247 2273 281
rect 2487 247 2503 281
rect 2537 247 2553 281
rect 2767 247 2783 281
rect 2817 247 2833 281
rect 3047 247 3063 281
rect 3097 247 3113 281
rect -61 188 -27 204
rect -61 -204 -27 -188
rect 27 188 61 204
rect 27 -204 61 -188
rect 219 188 253 204
rect 219 -204 253 -188
rect 307 188 341 204
rect 307 -204 341 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 587 188 621 204
rect 587 -204 621 -188
rect 779 188 813 204
rect 779 -204 813 -188
rect 867 188 901 204
rect 867 -204 901 -188
rect 1059 188 1093 204
rect 1059 -204 1093 -188
rect 1147 188 1181 204
rect 1147 -204 1181 -188
rect 1339 188 1373 204
rect 1339 -204 1373 -188
rect 1427 188 1461 204
rect 1427 -204 1461 -188
rect 1619 188 1653 204
rect 1619 -204 1653 -188
rect 1707 188 1741 204
rect 1707 -204 1741 -188
rect 1899 188 1933 204
rect 1899 -204 1933 -188
rect 1987 188 2021 204
rect 1987 -204 2021 -188
rect 2179 188 2213 204
rect 2179 -204 2213 -188
rect 2267 188 2301 204
rect 2267 -204 2301 -188
rect 2459 188 2493 204
rect 2459 -204 2493 -188
rect 2547 188 2581 204
rect 2547 -204 2581 -188
rect 2739 188 2773 204
rect 2739 -204 2773 -188
rect 2827 188 2861 204
rect 2827 -204 2861 -188
rect 3019 188 3053 204
rect 3019 -204 3053 -188
rect 3107 188 3141 204
rect 3107 -204 3141 -188
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect 247 -281 263 -247
rect 297 -281 313 -247
rect 527 -281 543 -247
rect 577 -281 593 -247
rect 807 -281 823 -247
rect 857 -281 873 -247
rect 1087 -281 1103 -247
rect 1137 -281 1153 -247
rect 1367 -281 1383 -247
rect 1417 -281 1433 -247
rect 1647 -281 1663 -247
rect 1697 -281 1713 -247
rect 1927 -281 1943 -247
rect 1977 -281 1993 -247
rect 2207 -281 2223 -247
rect 2257 -281 2273 -247
rect 2487 -281 2503 -247
rect 2537 -281 2553 -247
rect 2767 -281 2783 -247
rect 2817 -281 2833 -247
rect 3047 -281 3063 -247
rect 3097 -281 3113 -247
rect -33 -469 -17 -435
rect 17 -469 33 -435
rect 247 -469 263 -435
rect 297 -469 313 -435
rect 527 -469 543 -435
rect 577 -469 593 -435
rect 807 -469 823 -435
rect 857 -469 873 -435
rect 1087 -469 1103 -435
rect 1137 -469 1153 -435
rect 1367 -469 1383 -435
rect 1417 -469 1433 -435
rect 1647 -469 1663 -435
rect 1697 -469 1713 -435
rect 1927 -469 1943 -435
rect 1977 -469 1993 -435
rect 2207 -469 2223 -435
rect 2257 -469 2273 -435
rect 2487 -469 2503 -435
rect 2537 -469 2553 -435
rect 2767 -469 2783 -435
rect 2817 -469 2833 -435
rect 3047 -469 3063 -435
rect 3097 -469 3113 -435
rect -61 -528 -27 -512
rect -61 -920 -27 -904
rect 27 -528 61 -512
rect 27 -920 61 -904
rect 219 -528 253 -512
rect 219 -920 253 -904
rect 307 -528 341 -512
rect 307 -920 341 -904
rect 499 -528 533 -512
rect 499 -920 533 -904
rect 587 -528 621 -512
rect 587 -920 621 -904
rect 779 -528 813 -512
rect 779 -920 813 -904
rect 867 -528 901 -512
rect 867 -920 901 -904
rect 1059 -528 1093 -512
rect 1059 -920 1093 -904
rect 1147 -528 1181 -512
rect 1147 -920 1181 -904
rect 1339 -528 1373 -512
rect 1339 -920 1373 -904
rect 1427 -528 1461 -512
rect 1427 -920 1461 -904
rect 1619 -528 1653 -512
rect 1619 -920 1653 -904
rect 1707 -528 1741 -512
rect 1707 -920 1741 -904
rect 1899 -528 1933 -512
rect 1899 -920 1933 -904
rect 1987 -528 2021 -512
rect 1987 -920 2021 -904
rect 2179 -528 2213 -512
rect 2179 -920 2213 -904
rect 2267 -528 2301 -512
rect 2267 -920 2301 -904
rect 2459 -528 2493 -512
rect 2459 -920 2493 -904
rect 2547 -528 2581 -512
rect 2547 -920 2581 -904
rect 2739 -528 2773 -512
rect 2739 -920 2773 -904
rect 2827 -528 2861 -512
rect 2827 -920 2861 -904
rect 3019 -528 3053 -512
rect 3019 -920 3053 -904
rect 3107 -528 3141 -512
rect 3107 -920 3141 -904
rect -33 -997 -17 -963
rect 17 -997 33 -963
rect 247 -997 263 -963
rect 297 -997 313 -963
rect 527 -997 543 -963
rect 577 -997 593 -963
rect 807 -997 823 -963
rect 857 -997 873 -963
rect 1087 -997 1103 -963
rect 1137 -997 1153 -963
rect 1367 -997 1383 -963
rect 1417 -997 1433 -963
rect 1647 -997 1663 -963
rect 1697 -997 1713 -963
rect 1927 -997 1943 -963
rect 1977 -997 1993 -963
rect 2207 -997 2223 -963
rect 2257 -997 2273 -963
rect 2487 -997 2503 -963
rect 2537 -997 2553 -963
rect 2767 -997 2783 -963
rect 2817 -997 2833 -963
rect 3047 -997 3063 -963
rect 3097 -997 3113 -963
rect -496 -1702 -396 -1540
rect 3634 -1702 3734 -1540
rect -496 -2140 -396 -1978
rect 3634 -2140 3734 -1978
rect 246 -2571 262 -2537
rect 296 -2571 312 -2537
rect 526 -2571 542 -2537
rect 576 -2571 592 -2537
rect 806 -2571 822 -2537
rect 856 -2571 872 -2537
rect 1086 -2571 1102 -2537
rect 1136 -2571 1152 -2537
rect 1366 -2571 1382 -2537
rect 1416 -2571 1432 -2537
rect 1646 -2571 1662 -2537
rect 1696 -2571 1712 -2537
rect 1926 -2571 1942 -2537
rect 1976 -2571 1992 -2537
rect 2206 -2571 2222 -2537
rect 2256 -2571 2272 -2537
rect 2486 -2571 2502 -2537
rect 2536 -2571 2552 -2537
rect 2766 -2571 2782 -2537
rect 2816 -2571 2832 -2537
rect 218 -2621 252 -2605
rect 218 -3013 252 -2997
rect 306 -2621 340 -2605
rect 306 -3013 340 -2997
rect 498 -2621 532 -2605
rect 498 -3013 532 -2997
rect 586 -2621 620 -2605
rect 586 -3013 620 -2997
rect 778 -2621 812 -2605
rect 778 -3013 812 -2997
rect 866 -2621 900 -2605
rect 866 -3013 900 -2997
rect 1058 -2621 1092 -2605
rect 1058 -3013 1092 -2997
rect 1146 -2621 1180 -2605
rect 1146 -3013 1180 -2997
rect 1338 -2621 1372 -2605
rect 1338 -3013 1372 -2997
rect 1426 -2621 1460 -2605
rect 1426 -3013 1460 -2997
rect 1618 -2621 1652 -2605
rect 1618 -3013 1652 -2997
rect 1706 -2621 1740 -2605
rect 1706 -3013 1740 -2997
rect 1898 -2621 1932 -2605
rect 1898 -3013 1932 -2997
rect 1986 -2621 2020 -2605
rect 1986 -3013 2020 -2997
rect 2178 -2621 2212 -2605
rect 2178 -3013 2212 -2997
rect 2266 -2621 2300 -2605
rect 2266 -3013 2300 -2997
rect 2458 -2621 2492 -2605
rect 2458 -3013 2492 -2997
rect 2546 -2621 2580 -2605
rect 2546 -3013 2580 -2997
rect 2738 -2621 2772 -2605
rect 2738 -3013 2772 -2997
rect 2826 -2621 2860 -2605
rect 2826 -3013 2860 -2997
rect 246 -3081 262 -3047
rect 296 -3081 312 -3047
rect 526 -3081 542 -3047
rect 576 -3081 592 -3047
rect 806 -3081 822 -3047
rect 856 -3081 872 -3047
rect 1086 -3081 1102 -3047
rect 1136 -3081 1152 -3047
rect 1366 -3081 1382 -3047
rect 1416 -3081 1432 -3047
rect 1646 -3081 1662 -3047
rect 1696 -3081 1712 -3047
rect 1926 -3081 1942 -3047
rect 1976 -3081 1992 -3047
rect 2206 -3081 2222 -3047
rect 2256 -3081 2272 -3047
rect 2486 -3081 2502 -3047
rect 2536 -3081 2552 -3047
rect 2766 -3081 2782 -3047
rect 2816 -3081 2832 -3047
rect 246 -3391 262 -3357
rect 296 -3391 312 -3357
rect 526 -3391 542 -3357
rect 576 -3391 592 -3357
rect 806 -3391 822 -3357
rect 856 -3391 872 -3357
rect 1086 -3391 1102 -3357
rect 1136 -3391 1152 -3357
rect 1366 -3391 1382 -3357
rect 1416 -3391 1432 -3357
rect 1646 -3391 1662 -3357
rect 1696 -3391 1712 -3357
rect 1926 -3391 1942 -3357
rect 1976 -3391 1992 -3357
rect 2206 -3391 2222 -3357
rect 2256 -3391 2272 -3357
rect 2486 -3391 2502 -3357
rect 2536 -3391 2552 -3357
rect 2766 -3391 2782 -3357
rect 2816 -3391 2832 -3357
rect 218 -3441 252 -3425
rect 218 -3833 252 -3817
rect 306 -3441 340 -3425
rect 306 -3833 340 -3817
rect 498 -3441 532 -3425
rect 498 -3833 532 -3817
rect 586 -3441 620 -3425
rect 586 -3833 620 -3817
rect 778 -3441 812 -3425
rect 778 -3833 812 -3817
rect 866 -3441 900 -3425
rect 866 -3833 900 -3817
rect 1058 -3441 1092 -3425
rect 1058 -3833 1092 -3817
rect 1146 -3441 1180 -3425
rect 1146 -3833 1180 -3817
rect 1338 -3441 1372 -3425
rect 1338 -3833 1372 -3817
rect 1426 -3441 1460 -3425
rect 1426 -3833 1460 -3817
rect 1618 -3441 1652 -3425
rect 1618 -3833 1652 -3817
rect 1706 -3441 1740 -3425
rect 1706 -3833 1740 -3817
rect 1898 -3441 1932 -3425
rect 1898 -3833 1932 -3817
rect 1986 -3441 2020 -3425
rect 1986 -3833 2020 -3817
rect 2178 -3441 2212 -3425
rect 2178 -3833 2212 -3817
rect 2266 -3441 2300 -3425
rect 2266 -3833 2300 -3817
rect 2458 -3441 2492 -3425
rect 2458 -3833 2492 -3817
rect 2546 -3441 2580 -3425
rect 2546 -3833 2580 -3817
rect 2738 -3441 2772 -3425
rect 2738 -3833 2772 -3817
rect 2826 -3441 2860 -3425
rect 2826 -3833 2860 -3817
rect 246 -3901 262 -3867
rect 296 -3901 312 -3867
rect 526 -3901 542 -3867
rect 576 -3901 592 -3867
rect 806 -3901 822 -3867
rect 856 -3901 872 -3867
rect 1086 -3901 1102 -3867
rect 1136 -3901 1152 -3867
rect 1366 -3901 1382 -3867
rect 1416 -3901 1432 -3867
rect 1646 -3901 1662 -3867
rect 1696 -3901 1712 -3867
rect 1926 -3901 1942 -3867
rect 1976 -3901 1992 -3867
rect 2206 -3901 2222 -3867
rect 2256 -3901 2272 -3867
rect 2486 -3901 2502 -3867
rect 2536 -3901 2552 -3867
rect 2766 -3901 2782 -3867
rect 2816 -3901 2832 -3867
rect 1366 -4671 1382 -4637
rect 1416 -4671 1432 -4637
rect 1646 -4671 1662 -4637
rect 1696 -4671 1712 -4637
rect 1338 -4721 1372 -4705
rect 1338 -5113 1372 -5097
rect 1426 -4721 1460 -4705
rect 1426 -5113 1460 -5097
rect 1618 -4721 1652 -4705
rect 1618 -5113 1652 -5097
rect 1706 -4721 1740 -4705
rect 1706 -5113 1740 -5097
rect 1366 -5181 1382 -5147
rect 1416 -5181 1432 -5147
rect 1646 -5181 1662 -5147
rect 1696 -5181 1712 -5147
rect 1365 -5529 1381 -5495
rect 1415 -5529 1431 -5495
rect 1645 -5529 1661 -5495
rect 1695 -5529 1711 -5495
rect 1337 -5579 1371 -5563
rect 1337 -5971 1371 -5955
rect 1425 -5579 1459 -5563
rect 1425 -5971 1459 -5955
rect 1617 -5579 1651 -5563
rect 1617 -5971 1651 -5955
rect 1705 -5579 1739 -5563
rect 1705 -5971 1739 -5955
rect 246 -6474 262 -6440
rect 296 -6474 312 -6440
rect 526 -6474 542 -6440
rect 576 -6474 592 -6440
rect 806 -6474 822 -6440
rect 856 -6474 872 -6440
rect 1086 -6474 1102 -6440
rect 1136 -6474 1152 -6440
rect 1366 -6474 1382 -6440
rect 1416 -6474 1432 -6440
rect 1646 -6474 1662 -6440
rect 1696 -6474 1712 -6440
rect 1926 -6474 1942 -6440
rect 1976 -6474 1992 -6440
rect 2206 -6474 2222 -6440
rect 2256 -6474 2272 -6440
rect 2486 -6474 2502 -6440
rect 2536 -6474 2552 -6440
rect 2766 -6474 2782 -6440
rect 2816 -6474 2832 -6440
rect 218 -6524 252 -6508
rect 218 -6916 252 -6900
rect 306 -6524 340 -6508
rect 306 -6916 340 -6900
rect 498 -6524 532 -6508
rect 498 -6916 532 -6900
rect 586 -6524 620 -6508
rect 586 -6916 620 -6900
rect 778 -6524 812 -6508
rect 778 -6916 812 -6900
rect 866 -6524 900 -6508
rect 866 -6916 900 -6900
rect 1058 -6524 1092 -6508
rect 1058 -6916 1092 -6900
rect 1146 -6524 1180 -6508
rect 1146 -6916 1180 -6900
rect 1338 -6524 1372 -6508
rect 1338 -6916 1372 -6900
rect 1426 -6524 1460 -6508
rect 1426 -6916 1460 -6900
rect 1618 -6524 1652 -6508
rect 1618 -6916 1652 -6900
rect 1706 -6524 1740 -6508
rect 1706 -6916 1740 -6900
rect 1898 -6524 1932 -6508
rect 1898 -6916 1932 -6900
rect 1986 -6524 2020 -6508
rect 1986 -6916 2020 -6900
rect 2178 -6524 2212 -6508
rect 2178 -6916 2212 -6900
rect 2266 -6524 2300 -6508
rect 2266 -6916 2300 -6900
rect 2458 -6524 2492 -6508
rect 2458 -6916 2492 -6900
rect 2546 -6524 2580 -6508
rect 2546 -6916 2580 -6900
rect 2738 -6524 2772 -6508
rect 2738 -6916 2772 -6900
rect 2826 -6524 2860 -6508
rect 2826 -6916 2860 -6900
rect 218 -7222 252 -7206
rect 218 -7614 252 -7598
rect 306 -7222 340 -7206
rect 306 -7614 340 -7598
rect 498 -7222 532 -7206
rect 498 -7614 532 -7598
rect 586 -7222 620 -7206
rect 586 -7614 620 -7598
rect 778 -7222 812 -7206
rect 778 -7614 812 -7598
rect 866 -7222 900 -7206
rect 866 -7614 900 -7598
rect 1058 -7222 1092 -7206
rect 1058 -7614 1092 -7598
rect 1146 -7222 1180 -7206
rect 1146 -7614 1180 -7598
rect 1338 -7222 1372 -7206
rect 1338 -7614 1372 -7598
rect 1426 -7222 1460 -7206
rect 1426 -7614 1460 -7598
rect 1618 -7222 1652 -7206
rect 1618 -7614 1652 -7598
rect 1706 -7222 1740 -7206
rect 1706 -7614 1740 -7598
rect 1898 -7222 1932 -7206
rect 1898 -7614 1932 -7598
rect 1986 -7222 2020 -7206
rect 1986 -7614 2020 -7598
rect 2178 -7222 2212 -7206
rect 2178 -7614 2212 -7598
rect 2266 -7222 2300 -7206
rect 2266 -7614 2300 -7598
rect 2458 -7222 2492 -7206
rect 2458 -7614 2492 -7598
rect 2546 -7222 2580 -7206
rect 2546 -7614 2580 -7598
rect 2738 -7222 2772 -7206
rect 2738 -7614 2772 -7598
rect 2826 -7222 2860 -7206
rect 2826 -7614 2860 -7598
rect 246 -7682 262 -7648
rect 296 -7682 312 -7648
rect 526 -7682 542 -7648
rect 576 -7682 592 -7648
rect 806 -7682 822 -7648
rect 856 -7682 872 -7648
rect 1086 -7682 1102 -7648
rect 1136 -7682 1152 -7648
rect 1366 -7682 1382 -7648
rect 1416 -7682 1432 -7648
rect 1646 -7682 1662 -7648
rect 1696 -7682 1712 -7648
rect 1926 -7682 1942 -7648
rect 1976 -7682 1992 -7648
rect 2206 -7682 2222 -7648
rect 2256 -7682 2272 -7648
rect 2486 -7682 2502 -7648
rect 2536 -7682 2552 -7648
rect 2766 -7682 2782 -7648
rect 2816 -7682 2832 -7648
rect -496 -8594 -396 -8432
rect 3634 -8594 3734 -8432
<< viali >>
rect -396 1022 -334 1122
rect -334 1022 3572 1122
rect 3572 1022 3634 1122
rect -496 -1471 -396 891
rect -17 247 17 281
rect 263 247 297 281
rect 543 247 577 281
rect 823 247 857 281
rect 1103 247 1137 281
rect 1383 247 1417 281
rect 1663 247 1697 281
rect 1943 247 1977 281
rect 2223 247 2257 281
rect 2503 247 2537 281
rect 2783 247 2817 281
rect 3063 247 3097 281
rect -61 -188 -27 188
rect 27 -188 61 188
rect 219 -188 253 188
rect 307 -188 341 188
rect 499 -188 533 188
rect 587 -188 621 188
rect 779 -188 813 188
rect 867 -188 901 188
rect 1059 -188 1093 188
rect 1147 -188 1181 188
rect 1339 -188 1373 188
rect 1427 -188 1461 188
rect 1619 -188 1653 188
rect 1707 -188 1741 188
rect 1899 -188 1933 188
rect 1987 -188 2021 188
rect 2179 -188 2213 188
rect 2267 -188 2301 188
rect 2459 -188 2493 188
rect 2547 -188 2581 188
rect 2739 -188 2773 188
rect 2827 -188 2861 188
rect 3019 -188 3053 188
rect 3107 -188 3141 188
rect -17 -281 17 -247
rect 263 -281 297 -247
rect 543 -281 577 -247
rect 823 -281 857 -247
rect 1103 -281 1137 -247
rect 1383 -281 1417 -247
rect 1663 -281 1697 -247
rect 1943 -281 1977 -247
rect 2223 -281 2257 -247
rect 2503 -281 2537 -247
rect 2783 -281 2817 -247
rect 3063 -281 3097 -247
rect -17 -469 17 -435
rect 263 -469 297 -435
rect 543 -469 577 -435
rect 823 -469 857 -435
rect 1103 -469 1137 -435
rect 1383 -469 1417 -435
rect 1663 -469 1697 -435
rect 1943 -469 1977 -435
rect 2223 -469 2257 -435
rect 2503 -469 2537 -435
rect 2783 -469 2817 -435
rect 3063 -469 3097 -435
rect -61 -904 -27 -528
rect 27 -904 61 -528
rect 219 -904 253 -528
rect 307 -904 341 -528
rect 499 -904 533 -528
rect 587 -904 621 -528
rect 779 -904 813 -528
rect 867 -904 901 -528
rect 1059 -904 1093 -528
rect 1147 -904 1181 -528
rect 1339 -904 1373 -528
rect 1427 -904 1461 -528
rect 1619 -904 1653 -528
rect 1707 -904 1741 -528
rect 1899 -904 1933 -528
rect 1987 -904 2021 -528
rect 2179 -904 2213 -528
rect 2267 -904 2301 -528
rect 2459 -904 2493 -528
rect 2547 -904 2581 -528
rect 2739 -904 2773 -528
rect 2827 -904 2861 -528
rect 3019 -904 3053 -528
rect 3107 -904 3141 -528
rect -17 -997 17 -963
rect 263 -997 297 -963
rect 543 -997 577 -963
rect 823 -997 857 -963
rect 1103 -997 1137 -963
rect 1383 -997 1417 -963
rect 1663 -997 1697 -963
rect 1943 -997 1977 -963
rect 2223 -997 2257 -963
rect 2503 -997 2537 -963
rect 2783 -997 2817 -963
rect 3063 -997 3097 -963
rect 3634 -1471 3734 891
rect -396 -1702 -334 -1602
rect -334 -1702 3572 -1602
rect 3572 -1702 3634 -1602
rect -396 -2078 -334 -1978
rect -334 -2078 3572 -1978
rect 3572 -2078 3634 -1978
rect -496 -8162 -396 -2410
rect 262 -2571 296 -2537
rect 542 -2571 576 -2537
rect 822 -2571 856 -2537
rect 1102 -2571 1136 -2537
rect 1382 -2571 1416 -2537
rect 1662 -2571 1696 -2537
rect 1942 -2571 1976 -2537
rect 2222 -2571 2256 -2537
rect 2502 -2571 2536 -2537
rect 2782 -2571 2816 -2537
rect 218 -2997 252 -2621
rect 306 -2997 340 -2621
rect 498 -2997 532 -2621
rect 586 -2997 620 -2621
rect 778 -2997 812 -2621
rect 866 -2997 900 -2621
rect 1058 -2997 1092 -2621
rect 1146 -2997 1180 -2621
rect 1338 -2997 1372 -2621
rect 1426 -2997 1460 -2621
rect 1618 -2997 1652 -2621
rect 1706 -2997 1740 -2621
rect 1898 -2997 1932 -2621
rect 1986 -2997 2020 -2621
rect 2178 -2997 2212 -2621
rect 2266 -2997 2300 -2621
rect 2458 -2997 2492 -2621
rect 2546 -2997 2580 -2621
rect 2738 -2997 2772 -2621
rect 2826 -2997 2860 -2621
rect 262 -3081 296 -3047
rect 542 -3081 576 -3047
rect 822 -3081 856 -3047
rect 1102 -3081 1136 -3047
rect 1382 -3081 1416 -3047
rect 1662 -3081 1696 -3047
rect 1942 -3081 1976 -3047
rect 2222 -3081 2256 -3047
rect 2502 -3081 2536 -3047
rect 2782 -3081 2816 -3047
rect 262 -3391 296 -3357
rect 542 -3391 576 -3357
rect 822 -3391 856 -3357
rect 1102 -3391 1136 -3357
rect 1382 -3391 1416 -3357
rect 1662 -3391 1696 -3357
rect 1942 -3391 1976 -3357
rect 2222 -3391 2256 -3357
rect 2502 -3391 2536 -3357
rect 2782 -3391 2816 -3357
rect 218 -3817 252 -3441
rect 306 -3817 340 -3441
rect 498 -3817 532 -3441
rect 586 -3817 620 -3441
rect 778 -3817 812 -3441
rect 866 -3817 900 -3441
rect 1058 -3817 1092 -3441
rect 1146 -3817 1180 -3441
rect 1338 -3817 1372 -3441
rect 1426 -3817 1460 -3441
rect 1618 -3817 1652 -3441
rect 1706 -3817 1740 -3441
rect 1898 -3817 1932 -3441
rect 1986 -3817 2020 -3441
rect 2178 -3817 2212 -3441
rect 2266 -3817 2300 -3441
rect 2458 -3817 2492 -3441
rect 2546 -3817 2580 -3441
rect 2738 -3817 2772 -3441
rect 2826 -3817 2860 -3441
rect 262 -3901 296 -3867
rect 542 -3901 576 -3867
rect 822 -3901 856 -3867
rect 1102 -3901 1136 -3867
rect 1382 -3901 1416 -3867
rect 1662 -3901 1696 -3867
rect 1942 -3901 1976 -3867
rect 2222 -3901 2256 -3867
rect 2502 -3901 2536 -3867
rect 2782 -3901 2816 -3867
rect 1382 -4671 1416 -4637
rect 1662 -4671 1696 -4637
rect 1338 -5097 1372 -4721
rect 1426 -5097 1460 -4721
rect 1618 -5097 1652 -4721
rect 1706 -5097 1740 -4721
rect 1382 -5181 1416 -5147
rect 1662 -5181 1696 -5147
rect 1381 -5529 1415 -5495
rect 1661 -5529 1695 -5495
rect 1337 -5955 1371 -5579
rect 1425 -5955 1459 -5579
rect 1617 -5955 1651 -5579
rect 1705 -5955 1739 -5579
rect 262 -6474 296 -6440
rect 542 -6474 576 -6440
rect 822 -6474 856 -6440
rect 1102 -6474 1136 -6440
rect 1382 -6474 1416 -6440
rect 1662 -6474 1696 -6440
rect 1942 -6474 1976 -6440
rect 2222 -6474 2256 -6440
rect 2502 -6474 2536 -6440
rect 2782 -6474 2816 -6440
rect 218 -6900 252 -6524
rect 306 -6900 340 -6524
rect 498 -6900 532 -6524
rect 586 -6900 620 -6524
rect 778 -6900 812 -6524
rect 866 -6900 900 -6524
rect 1058 -6900 1092 -6524
rect 1146 -6900 1180 -6524
rect 1338 -6900 1372 -6524
rect 1426 -6900 1460 -6524
rect 1618 -6900 1652 -6524
rect 1706 -6900 1740 -6524
rect 1898 -6900 1932 -6524
rect 1986 -6900 2020 -6524
rect 2178 -6900 2212 -6524
rect 2266 -6900 2300 -6524
rect 2458 -6900 2492 -6524
rect 2546 -6900 2580 -6524
rect 2738 -6900 2772 -6524
rect 2826 -6900 2860 -6524
rect 218 -7598 252 -7222
rect 306 -7598 340 -7222
rect 498 -7598 532 -7222
rect 586 -7598 620 -7222
rect 778 -7598 812 -7222
rect 866 -7598 900 -7222
rect 1058 -7598 1092 -7222
rect 1146 -7598 1180 -7222
rect 1338 -7598 1372 -7222
rect 1426 -7598 1460 -7222
rect 1618 -7598 1652 -7222
rect 1706 -7598 1740 -7222
rect 1898 -7598 1932 -7222
rect 1986 -7598 2020 -7222
rect 2178 -7598 2212 -7222
rect 2266 -7598 2300 -7222
rect 2458 -7598 2492 -7222
rect 2546 -7598 2580 -7222
rect 2738 -7598 2772 -7222
rect 2826 -7598 2860 -7222
rect 262 -7682 296 -7648
rect 542 -7682 576 -7648
rect 822 -7682 856 -7648
rect 1102 -7682 1136 -7648
rect 1382 -7682 1416 -7648
rect 1662 -7682 1696 -7648
rect 1942 -7682 1976 -7648
rect 2222 -7682 2256 -7648
rect 2502 -7682 2536 -7648
rect 2782 -7682 2816 -7648
rect 3634 -8162 3734 -2410
rect -396 -8594 -334 -8494
rect -334 -8594 3572 -8494
rect 3572 -8594 3634 -8494
<< metal1 >>
rect -502 1122 3740 1128
rect -502 1022 -396 1122
rect 3634 1022 3740 1122
rect -502 1016 3740 1022
rect -502 891 -390 1016
rect -502 -1471 -496 891
rect -396 -1471 -390 891
rect 210 716 220 1016
rect 730 770 782 1016
rect 706 670 806 770
rect 3018 716 3028 1016
rect 3628 891 3740 1016
rect -110 492 -58 502
rect -110 200 -58 440
rect 170 492 222 502
rect -26 398 26 408
rect -26 336 26 346
rect -18 287 18 336
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect 170 200 222 440
rect 450 492 502 502
rect 254 398 306 408
rect 254 336 306 346
rect 262 287 298 336
rect 251 281 309 287
rect 251 247 263 281
rect 297 247 309 281
rect 251 241 309 247
rect 450 200 502 440
rect 730 492 782 670
rect 534 398 586 408
rect 534 336 586 346
rect 542 287 578 336
rect 531 281 589 287
rect 531 247 543 281
rect 577 247 589 281
rect 531 241 589 247
rect 730 200 782 440
rect 1010 492 1062 502
rect 814 398 866 408
rect 814 336 866 346
rect 822 287 858 336
rect 811 281 869 287
rect 811 247 823 281
rect 857 247 869 281
rect 811 241 869 247
rect 1010 200 1062 440
rect 1290 492 1342 502
rect 1094 398 1146 408
rect 1094 336 1146 346
rect 1102 287 1138 336
rect 1091 281 1149 287
rect 1091 247 1103 281
rect 1137 247 1149 281
rect 1091 241 1149 247
rect 1290 200 1342 440
rect 1570 492 1622 502
rect 1374 398 1426 408
rect 1374 336 1426 346
rect 1382 287 1418 336
rect 1371 281 1429 287
rect 1371 247 1383 281
rect 1417 247 1429 281
rect 1371 241 1429 247
rect 1570 200 1622 440
rect 1850 492 1902 502
rect 1654 398 1706 408
rect 1654 336 1706 346
rect 1662 287 1698 336
rect 1651 281 1709 287
rect 1651 247 1663 281
rect 1697 247 1709 281
rect 1651 241 1709 247
rect 1850 200 1902 440
rect 2130 492 2182 502
rect 1934 398 1986 408
rect 1934 336 1986 346
rect 1942 287 1978 336
rect 1931 281 1989 287
rect 1931 247 1943 281
rect 1977 247 1989 281
rect 1931 241 1989 247
rect 2130 200 2182 440
rect 2410 492 2462 502
rect 2214 398 2266 408
rect 2214 336 2266 346
rect 2222 287 2258 336
rect 2211 281 2269 287
rect 2211 247 2223 281
rect 2257 247 2269 281
rect 2211 241 2269 247
rect 2410 200 2462 440
rect 2690 492 2742 502
rect 2494 398 2546 408
rect 2494 336 2546 346
rect 2502 287 2538 336
rect 2491 281 2549 287
rect 2491 247 2503 281
rect 2537 247 2549 281
rect 2491 241 2549 247
rect 2690 200 2742 440
rect 2970 492 3022 502
rect 2774 398 2826 408
rect 2774 336 2826 346
rect 2782 287 2818 336
rect 2771 281 2829 287
rect 2771 247 2783 281
rect 2817 247 2829 281
rect 2771 241 2829 247
rect 2970 200 3022 440
rect 3051 282 3109 287
rect 3228 282 3238 290
rect 3051 281 3238 282
rect 3051 247 3063 281
rect 3097 247 3238 281
rect 3051 246 3238 247
rect 3051 241 3109 246
rect 3228 238 3238 246
rect 3290 238 3300 290
rect -110 188 -21 200
rect -110 -188 -61 188
rect -27 -188 -21 188
rect -110 -200 -21 -188
rect 21 188 67 200
rect 21 -188 27 188
rect 61 -30 67 188
rect 170 188 259 200
rect 61 -188 112 -30
rect 21 -200 112 -188
rect -110 -516 -58 -200
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
rect -18 -308 18 -287
rect 60 -330 112 -200
rect -18 -429 18 -408
rect -29 -435 29 -429
rect -29 -469 -17 -435
rect 17 -469 29 -435
rect -29 -475 29 -469
rect 60 -516 112 -382
rect -110 -528 -21 -516
rect -110 -684 -61 -528
rect -67 -904 -61 -684
rect -27 -904 -21 -528
rect -67 -916 -21 -904
rect 21 -528 112 -516
rect 21 -904 27 -528
rect 61 -904 112 -528
rect 170 -188 219 188
rect 253 -188 259 188
rect 170 -200 259 -188
rect 301 188 347 200
rect 301 -188 307 188
rect 341 -30 347 188
rect 450 188 539 200
rect 341 -188 392 -30
rect 301 -200 392 -188
rect 170 -516 222 -200
rect 251 -247 309 -241
rect 251 -281 263 -247
rect 297 -281 309 -247
rect 251 -287 309 -281
rect 262 -308 298 -287
rect 340 -330 392 -200
rect 262 -429 298 -408
rect 251 -435 309 -429
rect 251 -469 263 -435
rect 297 -469 309 -435
rect 251 -475 309 -469
rect 340 -516 392 -382
rect 170 -528 259 -516
rect 170 -684 219 -528
rect 21 -916 112 -904
rect 213 -904 219 -684
rect 253 -904 259 -528
rect 213 -916 259 -904
rect 301 -528 392 -516
rect 301 -904 307 -528
rect 341 -682 392 -528
rect 450 -188 499 188
rect 533 -188 539 188
rect 450 -200 539 -188
rect 581 188 627 200
rect 581 -188 587 188
rect 621 -30 627 188
rect 730 188 819 200
rect 621 -188 672 -30
rect 581 -200 672 -188
rect 450 -516 502 -200
rect 531 -247 589 -241
rect 531 -281 543 -247
rect 577 -281 589 -247
rect 531 -287 589 -281
rect 542 -308 578 -287
rect 620 -330 672 -200
rect 542 -429 578 -408
rect 531 -435 589 -429
rect 531 -469 543 -435
rect 577 -469 589 -435
rect 531 -475 589 -469
rect 620 -516 672 -382
rect 450 -528 539 -516
rect 341 -904 347 -682
rect 450 -684 499 -528
rect 301 -916 347 -904
rect 493 -904 499 -684
rect 533 -904 539 -528
rect 493 -916 539 -904
rect 581 -528 672 -516
rect 581 -904 587 -528
rect 621 -682 672 -528
rect 730 -188 779 188
rect 813 -188 819 188
rect 730 -200 819 -188
rect 861 188 907 200
rect 861 -188 867 188
rect 901 -30 907 188
rect 1010 188 1099 200
rect 901 -188 952 -30
rect 861 -200 952 -188
rect 730 -516 782 -200
rect 811 -247 869 -241
rect 811 -281 823 -247
rect 857 -281 869 -247
rect 811 -287 869 -281
rect 822 -308 858 -287
rect 900 -330 952 -200
rect 822 -429 858 -408
rect 811 -435 869 -429
rect 811 -469 823 -435
rect 857 -469 869 -435
rect 811 -475 869 -469
rect 900 -516 952 -382
rect 730 -528 819 -516
rect 621 -904 627 -682
rect 730 -684 779 -528
rect 581 -916 627 -904
rect 773 -904 779 -684
rect 813 -904 819 -528
rect 773 -916 819 -904
rect 861 -528 952 -516
rect 861 -904 867 -528
rect 901 -682 952 -528
rect 1010 -188 1059 188
rect 1093 -188 1099 188
rect 1010 -200 1099 -188
rect 1141 188 1187 200
rect 1141 -188 1147 188
rect 1181 -30 1187 188
rect 1290 188 1379 200
rect 1181 -188 1232 -30
rect 1141 -200 1232 -188
rect 1010 -516 1062 -200
rect 1091 -247 1149 -241
rect 1091 -281 1103 -247
rect 1137 -281 1149 -247
rect 1091 -287 1149 -281
rect 1102 -308 1138 -287
rect 1180 -330 1232 -200
rect 1102 -429 1138 -408
rect 1091 -435 1149 -429
rect 1091 -469 1103 -435
rect 1137 -469 1149 -435
rect 1091 -475 1149 -469
rect 1180 -516 1232 -382
rect 1010 -528 1099 -516
rect 901 -904 907 -682
rect 1010 -684 1059 -528
rect 861 -916 907 -904
rect 1053 -904 1059 -684
rect 1093 -904 1099 -528
rect 1053 -916 1099 -904
rect 1141 -528 1232 -516
rect 1141 -904 1147 -528
rect 1181 -682 1232 -528
rect 1290 -188 1339 188
rect 1373 -188 1379 188
rect 1290 -200 1379 -188
rect 1421 188 1467 200
rect 1421 -188 1427 188
rect 1461 -30 1467 188
rect 1570 188 1659 200
rect 1461 -188 1512 -30
rect 1421 -200 1512 -188
rect 1290 -516 1342 -200
rect 1371 -247 1429 -241
rect 1371 -281 1383 -247
rect 1417 -281 1429 -247
rect 1371 -287 1429 -281
rect 1382 -308 1418 -287
rect 1460 -330 1512 -200
rect 1382 -429 1418 -408
rect 1371 -435 1429 -429
rect 1371 -469 1383 -435
rect 1417 -469 1429 -435
rect 1371 -475 1429 -469
rect 1460 -516 1512 -382
rect 1290 -528 1379 -516
rect 1181 -904 1187 -682
rect 1290 -684 1339 -528
rect 1141 -916 1187 -904
rect 1333 -904 1339 -684
rect 1373 -904 1379 -528
rect 1333 -916 1379 -904
rect 1421 -528 1512 -516
rect 1421 -904 1427 -528
rect 1461 -682 1512 -528
rect 1570 -188 1619 188
rect 1653 -188 1659 188
rect 1570 -200 1659 -188
rect 1701 188 1747 200
rect 1701 -188 1707 188
rect 1741 -30 1747 188
rect 1850 188 1939 200
rect 1741 -188 1792 -30
rect 1701 -200 1792 -188
rect 1570 -516 1622 -200
rect 1651 -247 1709 -241
rect 1651 -281 1663 -247
rect 1697 -281 1709 -247
rect 1651 -287 1709 -281
rect 1662 -308 1698 -287
rect 1740 -330 1792 -200
rect 1662 -429 1698 -408
rect 1651 -435 1709 -429
rect 1651 -469 1663 -435
rect 1697 -469 1709 -435
rect 1651 -475 1709 -469
rect 1740 -516 1792 -382
rect 1570 -528 1659 -516
rect 1461 -904 1467 -682
rect 1570 -684 1619 -528
rect 1421 -916 1467 -904
rect 1613 -904 1619 -684
rect 1653 -904 1659 -528
rect 1613 -916 1659 -904
rect 1701 -528 1792 -516
rect 1701 -904 1707 -528
rect 1741 -682 1792 -528
rect 1850 -188 1899 188
rect 1933 -188 1939 188
rect 1850 -200 1939 -188
rect 1981 188 2027 200
rect 1981 -188 1987 188
rect 2021 -30 2027 188
rect 2130 188 2219 200
rect 2021 -188 2072 -30
rect 1981 -200 2072 -188
rect 1850 -516 1902 -200
rect 1931 -247 1989 -241
rect 1931 -281 1943 -247
rect 1977 -281 1989 -247
rect 1931 -287 1989 -281
rect 1942 -308 1978 -287
rect 2020 -330 2072 -200
rect 1942 -429 1978 -408
rect 1931 -435 1989 -429
rect 1931 -469 1943 -435
rect 1977 -469 1989 -435
rect 1931 -475 1989 -469
rect 2020 -516 2072 -382
rect 1850 -528 1939 -516
rect 1741 -904 1747 -682
rect 1850 -684 1899 -528
rect 1701 -916 1747 -904
rect 1893 -904 1899 -684
rect 1933 -904 1939 -528
rect 1893 -916 1939 -904
rect 1981 -528 2072 -516
rect 1981 -904 1987 -528
rect 2021 -682 2072 -528
rect 2130 -188 2179 188
rect 2213 -188 2219 188
rect 2130 -200 2219 -188
rect 2261 188 2307 200
rect 2261 -188 2267 188
rect 2301 -30 2307 188
rect 2410 188 2499 200
rect 2301 -188 2352 -30
rect 2261 -200 2352 -188
rect 2130 -516 2182 -200
rect 2211 -247 2269 -241
rect 2211 -281 2223 -247
rect 2257 -281 2269 -247
rect 2211 -287 2269 -281
rect 2222 -308 2258 -287
rect 2300 -330 2352 -200
rect 2222 -429 2258 -408
rect 2211 -435 2269 -429
rect 2211 -469 2223 -435
rect 2257 -469 2269 -435
rect 2211 -475 2269 -469
rect 2300 -516 2352 -382
rect 2130 -528 2219 -516
rect 2021 -904 2027 -682
rect 2130 -684 2179 -528
rect 1981 -916 2027 -904
rect 2173 -904 2179 -684
rect 2213 -904 2219 -528
rect 2173 -916 2219 -904
rect 2261 -528 2352 -516
rect 2261 -904 2267 -528
rect 2301 -682 2352 -528
rect 2410 -188 2459 188
rect 2493 -188 2499 188
rect 2410 -200 2499 -188
rect 2541 188 2587 200
rect 2541 -188 2547 188
rect 2581 -30 2587 188
rect 2690 188 2779 200
rect 2581 -188 2632 -30
rect 2541 -200 2632 -188
rect 2410 -516 2462 -200
rect 2491 -247 2549 -241
rect 2491 -281 2503 -247
rect 2537 -281 2549 -247
rect 2491 -287 2549 -281
rect 2502 -308 2538 -287
rect 2580 -330 2632 -200
rect 2502 -429 2538 -408
rect 2491 -435 2549 -429
rect 2491 -469 2503 -435
rect 2537 -469 2549 -435
rect 2491 -475 2549 -469
rect 2580 -516 2632 -382
rect 2410 -528 2499 -516
rect 2301 -904 2307 -682
rect 2410 -684 2459 -528
rect 2261 -916 2307 -904
rect 2453 -904 2459 -684
rect 2493 -904 2499 -528
rect 2453 -916 2499 -904
rect 2541 -528 2632 -516
rect 2541 -904 2547 -528
rect 2581 -682 2632 -528
rect 2690 -188 2739 188
rect 2773 -188 2779 188
rect 2690 -200 2779 -188
rect 2821 188 2867 200
rect 2821 -188 2827 188
rect 2861 -30 2867 188
rect 2970 188 3059 200
rect 2861 -188 2912 -30
rect 2821 -200 2912 -188
rect 2690 -516 2742 -200
rect 2771 -247 2829 -241
rect 2771 -281 2783 -247
rect 2817 -281 2829 -247
rect 2771 -287 2829 -281
rect 2782 -308 2818 -287
rect 2860 -330 2912 -200
rect 2782 -429 2818 -408
rect 2771 -435 2829 -429
rect 2771 -469 2783 -435
rect 2817 -469 2829 -435
rect 2771 -475 2829 -469
rect 2860 -516 2912 -382
rect 2690 -528 2779 -516
rect 2581 -904 2587 -682
rect 2690 -684 2739 -528
rect 2541 -916 2587 -904
rect 2733 -904 2739 -684
rect 2773 -904 2779 -528
rect 2733 -916 2779 -904
rect 2821 -528 2912 -516
rect 2821 -904 2827 -528
rect 2861 -682 2912 -528
rect 2970 -188 3019 188
rect 3053 -188 3059 188
rect 2970 -200 3059 -188
rect 3101 188 3147 200
rect 3101 -188 3107 188
rect 3141 -30 3147 188
rect 3141 -188 3192 -30
rect 3101 -200 3192 -188
rect 2970 -516 3022 -200
rect 3051 -247 3109 -241
rect 3051 -281 3063 -247
rect 3097 -281 3109 -247
rect 3051 -287 3109 -281
rect 3062 -308 3098 -287
rect 3140 -330 3192 -200
rect 3062 -429 3098 -408
rect 3051 -435 3109 -429
rect 3051 -469 3063 -435
rect 3097 -469 3109 -435
rect 3051 -475 3109 -469
rect 3140 -516 3192 -382
rect 2970 -528 3059 -516
rect 2861 -904 2867 -682
rect 2970 -684 3019 -528
rect 2821 -916 2867 -904
rect 3013 -904 3019 -684
rect 3053 -904 3059 -528
rect 3013 -916 3059 -904
rect 3101 -528 3192 -516
rect 3101 -904 3107 -528
rect 3141 -904 3192 -528
rect 3101 -916 3192 -904
rect -29 -963 29 -957
rect -29 -997 -17 -963
rect 17 -997 29 -963
rect -29 -1003 29 -997
rect -18 -1052 18 -1003
rect -26 -1062 26 -1052
rect -26 -1124 26 -1114
rect 60 -1300 112 -916
rect 251 -963 309 -957
rect 251 -997 263 -963
rect 297 -997 309 -963
rect 251 -1003 309 -997
rect 531 -963 589 -957
rect 531 -997 543 -963
rect 577 -997 589 -963
rect 531 -1003 589 -997
rect 811 -963 869 -957
rect 811 -997 823 -963
rect 857 -997 869 -963
rect 811 -1003 869 -997
rect 1091 -963 1149 -957
rect 1091 -997 1103 -963
rect 1137 -997 1149 -963
rect 1091 -1003 1149 -997
rect 1371 -963 1429 -957
rect 1371 -997 1383 -963
rect 1417 -997 1429 -963
rect 1371 -1003 1429 -997
rect 1651 -963 1709 -957
rect 1651 -997 1663 -963
rect 1697 -997 1709 -963
rect 1651 -1003 1709 -997
rect 1931 -963 1989 -957
rect 1931 -997 1943 -963
rect 1977 -997 1989 -963
rect 1931 -1003 1989 -997
rect 2211 -963 2269 -957
rect 2211 -997 2223 -963
rect 2257 -997 2269 -963
rect 2211 -1003 2269 -997
rect 2491 -963 2549 -957
rect 2491 -997 2503 -963
rect 2537 -997 2549 -963
rect 2491 -1003 2549 -997
rect 2771 -963 2829 -957
rect 2771 -997 2783 -963
rect 2817 -997 2829 -963
rect 2771 -1003 2829 -997
rect 3051 -963 3109 -957
rect 3051 -997 3063 -963
rect 3097 -997 3109 -963
rect 3051 -1003 3109 -997
rect 262 -1052 298 -1003
rect 542 -1052 578 -1003
rect 822 -1052 858 -1003
rect 1102 -1052 1138 -1003
rect 254 -1062 306 -1052
rect 254 -1124 306 -1114
rect 534 -1062 586 -1052
rect 534 -1124 586 -1114
rect 814 -1062 866 -1052
rect 814 -1124 866 -1114
rect 1094 -1062 1146 -1052
rect 1094 -1124 1146 -1114
rect 1382 -1168 1418 -1003
rect 1662 -1168 1698 -1003
rect 1942 -1052 1978 -1003
rect 2222 -1052 2258 -1003
rect 2502 -1052 2538 -1003
rect 2782 -1052 2818 -1003
rect 3062 -1052 3098 -1003
rect 1934 -1062 1986 -1052
rect 1934 -1124 1986 -1114
rect 2214 -1062 2266 -1052
rect 2214 -1124 2266 -1114
rect 2494 -1062 2546 -1052
rect 2494 -1124 2546 -1114
rect 2774 -1062 2826 -1052
rect 2774 -1124 2826 -1114
rect 3054 -1062 3106 -1052
rect 3054 -1124 3106 -1114
rect 1374 -1178 1426 -1168
rect 1374 -1240 1426 -1230
rect 1654 -1178 1706 -1168
rect 1654 -1240 1706 -1230
rect 34 -1400 134 -1300
rect -502 -1596 -390 -1471
rect 66 -1472 102 -1400
rect 404 -1472 414 -1462
rect 66 -1508 414 -1472
rect 404 -1514 414 -1508
rect 466 -1472 476 -1462
rect 1662 -1472 1698 -1240
rect 2368 -1372 2468 -1348
rect 3140 -1372 3192 -916
rect 2368 -1424 2478 -1372
rect 2530 -1424 3192 -1372
rect 2368 -1448 2468 -1424
rect 466 -1508 1698 -1472
rect 3628 -1471 3634 891
rect 3734 -1471 3740 891
rect 466 -1514 476 -1508
rect 3628 -1596 3740 -1471
rect -502 -1602 3740 -1596
rect -502 -1702 -396 -1602
rect 3634 -1702 3740 -1602
rect -502 -1708 3740 -1702
rect 2906 -1862 2916 -1810
rect 2968 -1816 2978 -1810
rect 3274 -1816 3374 -1792
rect 2968 -1854 3374 -1816
rect 2968 -1862 2978 -1854
rect 3274 -1892 3374 -1854
rect -502 -1978 3740 -1972
rect -502 -2078 -396 -1978
rect 3634 -2078 3740 -1978
rect -502 -2084 3740 -2078
rect -502 -2410 -390 -2084
rect 900 -2142 952 -2132
rect 900 -2204 952 -2194
rect 2774 -2134 2826 -2124
rect 2774 -2196 2826 -2186
rect 330 -2222 382 -2212
rect 330 -2284 382 -2274
rect 610 -2222 662 -2212
rect 610 -2284 662 -2274
rect 178 -2322 230 -2312
rect 178 -2384 230 -2374
rect -502 -8162 -496 -2410
rect -396 -8162 -390 -2410
rect 186 -2609 222 -2384
rect 254 -2422 306 -2412
rect 254 -2484 306 -2474
rect 262 -2531 298 -2484
rect 250 -2537 308 -2531
rect 250 -2571 262 -2537
rect 296 -2571 308 -2537
rect 250 -2577 308 -2571
rect 338 -2609 374 -2284
rect 458 -2322 510 -2312
rect 458 -2384 510 -2374
rect 186 -2621 258 -2609
rect 186 -2670 218 -2621
rect 212 -2997 218 -2670
rect 252 -2997 258 -2621
rect 212 -3009 258 -2997
rect 300 -2621 374 -2609
rect 300 -2997 306 -2621
rect 340 -2670 374 -2621
rect 466 -2609 502 -2384
rect 534 -2422 586 -2412
rect 534 -2484 586 -2474
rect 542 -2531 578 -2484
rect 530 -2537 588 -2531
rect 530 -2571 542 -2537
rect 576 -2571 588 -2537
rect 530 -2577 588 -2571
rect 618 -2609 654 -2284
rect 814 -2422 866 -2412
rect 814 -2484 866 -2474
rect 822 -2531 858 -2484
rect 810 -2537 868 -2531
rect 810 -2571 822 -2537
rect 856 -2571 868 -2537
rect 810 -2577 868 -2571
rect 900 -2609 936 -2204
rect 1450 -2222 1502 -2212
rect 1450 -2284 1502 -2274
rect 1730 -2222 1782 -2212
rect 1730 -2284 1782 -2274
rect 2570 -2222 2622 -2212
rect 2570 -2284 2622 -2274
rect 1298 -2322 1350 -2312
rect 1298 -2384 1350 -2374
rect 1094 -2422 1146 -2412
rect 1094 -2484 1146 -2474
rect 1102 -2531 1138 -2484
rect 1090 -2537 1148 -2531
rect 1090 -2571 1102 -2537
rect 1136 -2571 1148 -2537
rect 1090 -2577 1148 -2571
rect 1306 -2609 1342 -2384
rect 1374 -2422 1426 -2412
rect 1374 -2484 1426 -2474
rect 1382 -2531 1418 -2484
rect 1370 -2537 1428 -2531
rect 1370 -2571 1382 -2537
rect 1416 -2571 1428 -2537
rect 1370 -2577 1428 -2571
rect 1458 -2609 1494 -2284
rect 1578 -2322 1630 -2312
rect 1578 -2384 1630 -2374
rect 466 -2621 538 -2609
rect 466 -2670 498 -2621
rect 340 -2997 346 -2670
rect 300 -3009 346 -2997
rect 492 -2997 498 -2670
rect 532 -2997 538 -2621
rect 492 -3009 538 -2997
rect 580 -2621 654 -2609
rect 580 -2997 586 -2621
rect 620 -2670 654 -2621
rect 772 -2621 818 -2609
rect 620 -2997 626 -2670
rect 772 -2950 778 -2621
rect 580 -3009 626 -2997
rect 746 -2997 778 -2950
rect 812 -2997 818 -2621
rect 746 -3009 818 -2997
rect 860 -2621 936 -2609
rect 860 -2997 866 -2621
rect 900 -2997 936 -2621
rect 1052 -2621 1098 -2609
rect 1052 -2950 1058 -2621
rect 860 -3009 936 -2997
rect 250 -3047 308 -3041
rect 250 -3081 262 -3047
rect 296 -3081 308 -3047
rect 250 -3087 308 -3081
rect 530 -3047 588 -3041
rect 530 -3081 542 -3047
rect 576 -3081 588 -3047
rect 530 -3087 588 -3081
rect 262 -3108 298 -3087
rect 542 -3108 578 -3087
rect 746 -3132 782 -3009
rect 810 -3047 868 -3041
rect 810 -3081 822 -3047
rect 856 -3081 868 -3047
rect 810 -3087 868 -3081
rect 898 -3054 936 -3009
rect 1026 -2997 1058 -2950
rect 1092 -2997 1098 -2621
rect 1026 -3009 1098 -2997
rect 1140 -2621 1186 -2609
rect 1140 -2997 1146 -2621
rect 1180 -2950 1186 -2621
rect 1306 -2621 1378 -2609
rect 1306 -2670 1338 -2621
rect 1180 -2997 1214 -2950
rect 1140 -3009 1214 -2997
rect 1332 -2997 1338 -2670
rect 1372 -2997 1378 -2621
rect 1332 -3009 1378 -2997
rect 1420 -2621 1494 -2609
rect 1420 -2997 1426 -2621
rect 1460 -2670 1494 -2621
rect 1586 -2609 1622 -2384
rect 1654 -2422 1706 -2412
rect 1654 -2484 1706 -2474
rect 1662 -2531 1698 -2484
rect 1650 -2537 1708 -2531
rect 1650 -2571 1662 -2537
rect 1696 -2571 1708 -2537
rect 1650 -2577 1708 -2571
rect 1738 -2609 1774 -2284
rect 2418 -2322 2470 -2312
rect 2418 -2384 2470 -2374
rect 1934 -2422 1986 -2412
rect 1934 -2484 1986 -2474
rect 2214 -2422 2266 -2412
rect 2214 -2484 2266 -2474
rect 1942 -2531 1978 -2484
rect 2222 -2531 2258 -2484
rect 1930 -2537 1988 -2531
rect 1930 -2571 1942 -2537
rect 1976 -2571 1988 -2537
rect 1930 -2577 1988 -2571
rect 2210 -2537 2268 -2531
rect 2210 -2571 2222 -2537
rect 2256 -2571 2268 -2537
rect 2210 -2577 2268 -2571
rect 2426 -2609 2462 -2384
rect 2494 -2422 2546 -2412
rect 2494 -2484 2546 -2474
rect 2502 -2531 2538 -2484
rect 2490 -2537 2548 -2531
rect 2490 -2571 2502 -2537
rect 2536 -2571 2548 -2537
rect 2490 -2577 2548 -2571
rect 2578 -2609 2614 -2284
rect 2698 -2322 2750 -2312
rect 2698 -2384 2750 -2374
rect 1586 -2621 1658 -2609
rect 1586 -2670 1618 -2621
rect 1460 -2997 1466 -2670
rect 1420 -3009 1466 -2997
rect 1612 -2997 1618 -2670
rect 1652 -2997 1658 -2621
rect 1612 -3009 1658 -2997
rect 1700 -2621 1774 -2609
rect 1700 -2997 1706 -2621
rect 1740 -2670 1774 -2621
rect 1892 -2621 1938 -2609
rect 1740 -2997 1746 -2670
rect 1892 -2950 1898 -2621
rect 1700 -3009 1746 -2997
rect 1866 -2997 1898 -2950
rect 1932 -2997 1938 -2621
rect 1866 -3009 1938 -2997
rect 1980 -2621 2026 -2609
rect 1980 -2997 1986 -2621
rect 2020 -2950 2026 -2621
rect 2172 -2621 2218 -2609
rect 2172 -2950 2178 -2621
rect 2020 -2997 2054 -2950
rect 1980 -3009 2054 -2997
rect 822 -3108 858 -3087
rect 178 -3146 230 -3136
rect 178 -3208 230 -3198
rect 458 -3146 510 -3136
rect 458 -3208 510 -3198
rect 738 -3142 790 -3132
rect 738 -3204 790 -3194
rect 186 -3429 222 -3208
rect 330 -3246 382 -3236
rect 330 -3308 382 -3298
rect 262 -3351 298 -3332
rect 250 -3357 308 -3351
rect 250 -3391 262 -3357
rect 296 -3391 308 -3357
rect 250 -3397 308 -3391
rect 338 -3429 374 -3308
rect 186 -3441 258 -3429
rect 186 -3488 218 -3441
rect 212 -3817 218 -3488
rect 252 -3817 258 -3441
rect 212 -3829 258 -3817
rect 300 -3441 374 -3429
rect 300 -3817 306 -3441
rect 340 -3490 374 -3441
rect 466 -3429 502 -3208
rect 898 -3236 934 -3054
rect 1026 -3132 1062 -3009
rect 1090 -3047 1148 -3041
rect 1090 -3081 1102 -3047
rect 1136 -3081 1148 -3047
rect 1090 -3087 1148 -3081
rect 1102 -3108 1138 -3087
rect 1018 -3142 1070 -3132
rect 1018 -3204 1070 -3194
rect 1178 -3236 1214 -3009
rect 1370 -3047 1428 -3041
rect 1370 -3081 1382 -3047
rect 1416 -3081 1428 -3047
rect 1370 -3087 1428 -3081
rect 1650 -3047 1708 -3041
rect 1650 -3081 1662 -3047
rect 1696 -3081 1708 -3047
rect 1650 -3087 1708 -3081
rect 1382 -3108 1418 -3087
rect 1662 -3108 1698 -3087
rect 1866 -3132 1902 -3009
rect 1930 -3047 1988 -3041
rect 1930 -3081 1942 -3047
rect 1976 -3081 1988 -3047
rect 1930 -3087 1988 -3081
rect 1942 -3108 1978 -3087
rect 1298 -3146 1350 -3136
rect 1298 -3208 1350 -3198
rect 1578 -3146 1630 -3136
rect 1578 -3208 1630 -3198
rect 1858 -3142 1910 -3132
rect 1858 -3204 1910 -3194
rect 610 -3246 662 -3236
rect 610 -3308 662 -3298
rect 890 -3246 942 -3236
rect 890 -3308 942 -3298
rect 1170 -3246 1222 -3236
rect 1170 -3308 1222 -3298
rect 542 -3351 578 -3332
rect 530 -3357 588 -3351
rect 530 -3391 542 -3357
rect 576 -3391 588 -3357
rect 530 -3397 588 -3391
rect 618 -3429 654 -3308
rect 822 -3351 858 -3332
rect 1102 -3351 1138 -3332
rect 810 -3357 868 -3351
rect 810 -3391 822 -3357
rect 856 -3391 868 -3357
rect 810 -3397 868 -3391
rect 1090 -3357 1148 -3351
rect 1090 -3391 1102 -3357
rect 1136 -3391 1148 -3357
rect 1090 -3397 1148 -3391
rect 1306 -3429 1342 -3208
rect 1450 -3246 1502 -3236
rect 1450 -3308 1502 -3298
rect 1382 -3351 1418 -3332
rect 1370 -3357 1428 -3351
rect 1370 -3391 1382 -3357
rect 1416 -3391 1428 -3357
rect 1370 -3397 1428 -3391
rect 1458 -3429 1494 -3308
rect 466 -3441 538 -3429
rect 466 -3490 498 -3441
rect 340 -3817 346 -3490
rect 300 -3829 346 -3817
rect 492 -3817 498 -3490
rect 532 -3817 538 -3441
rect 492 -3829 538 -3817
rect 580 -3441 654 -3429
rect 580 -3817 586 -3441
rect 620 -3490 654 -3441
rect 772 -3441 818 -3429
rect 620 -3817 626 -3490
rect 772 -3770 778 -3441
rect 580 -3829 626 -3817
rect 746 -3817 778 -3770
rect 812 -3817 818 -3441
rect 746 -3829 818 -3817
rect 860 -3441 906 -3429
rect 860 -3817 866 -3441
rect 900 -3770 906 -3441
rect 1052 -3441 1098 -3429
rect 1052 -3770 1058 -3441
rect 900 -3817 934 -3770
rect 860 -3829 934 -3817
rect 250 -3867 308 -3861
rect 250 -3901 262 -3867
rect 296 -3901 308 -3867
rect 250 -3907 308 -3901
rect 530 -3867 588 -3861
rect 530 -3901 542 -3867
rect 576 -3901 588 -3867
rect 530 -3907 588 -3901
rect 262 -3956 298 -3907
rect 542 -3956 578 -3907
rect 254 -3966 306 -3956
rect 254 -4028 306 -4018
rect 534 -3966 586 -3956
rect 534 -4028 586 -4018
rect 746 -4156 782 -3829
rect 810 -3867 868 -3861
rect 810 -3901 822 -3867
rect 856 -3901 868 -3867
rect 810 -3907 868 -3901
rect 822 -3956 858 -3907
rect 814 -3966 866 -3956
rect 814 -4028 866 -4018
rect 898 -4056 934 -3829
rect 1026 -3817 1058 -3770
rect 1092 -3817 1098 -3441
rect 1026 -3829 1098 -3817
rect 1140 -3441 1186 -3429
rect 1140 -3817 1146 -3441
rect 1180 -3770 1186 -3441
rect 1306 -3441 1378 -3429
rect 1306 -3490 1338 -3441
rect 1180 -3817 1214 -3770
rect 1140 -3829 1214 -3817
rect 1332 -3817 1338 -3490
rect 1372 -3817 1378 -3441
rect 1332 -3829 1378 -3817
rect 1420 -3441 1494 -3429
rect 1420 -3817 1426 -3441
rect 1460 -3490 1494 -3441
rect 1586 -3429 1622 -3208
rect 2018 -3236 2054 -3009
rect 2146 -2997 2178 -2950
rect 2212 -2997 2218 -2621
rect 2146 -3009 2218 -2997
rect 2260 -2621 2306 -2609
rect 2260 -2997 2266 -2621
rect 2300 -2950 2306 -2621
rect 2426 -2621 2498 -2609
rect 2426 -2670 2458 -2621
rect 2300 -2997 2334 -2950
rect 2260 -3009 2334 -2997
rect 2452 -2997 2458 -2670
rect 2492 -2997 2498 -2621
rect 2452 -3009 2498 -2997
rect 2540 -2621 2614 -2609
rect 2540 -2997 2546 -2621
rect 2580 -2670 2614 -2621
rect 2706 -2609 2742 -2384
rect 2782 -2412 2818 -2196
rect 2850 -2222 2902 -2212
rect 2850 -2284 2902 -2274
rect 2774 -2422 2826 -2412
rect 2774 -2484 2826 -2474
rect 2782 -2531 2818 -2484
rect 2770 -2537 2828 -2531
rect 2770 -2571 2782 -2537
rect 2816 -2571 2828 -2537
rect 2770 -2577 2828 -2571
rect 2858 -2609 2894 -2284
rect 2706 -2621 2778 -2609
rect 2706 -2670 2738 -2621
rect 2580 -2997 2586 -2670
rect 2540 -3009 2586 -2997
rect 2732 -2997 2738 -2670
rect 2772 -2997 2778 -2621
rect 2732 -3009 2778 -2997
rect 2820 -2621 2894 -2609
rect 2820 -2997 2826 -2621
rect 2860 -2670 2894 -2621
rect 3628 -2410 3740 -2084
rect 2860 -2997 2866 -2670
rect 2820 -3009 2866 -2997
rect 2146 -3132 2182 -3009
rect 2210 -3047 2268 -3041
rect 2210 -3081 2222 -3047
rect 2256 -3081 2268 -3047
rect 2210 -3087 2268 -3081
rect 2222 -3108 2258 -3087
rect 2138 -3142 2190 -3132
rect 2138 -3204 2190 -3194
rect 2298 -3236 2334 -3009
rect 2490 -3047 2548 -3041
rect 2490 -3081 2502 -3047
rect 2536 -3081 2548 -3047
rect 2490 -3087 2548 -3081
rect 2770 -3047 2828 -3041
rect 2770 -3081 2782 -3047
rect 2816 -3081 2828 -3047
rect 2770 -3087 2828 -3081
rect 2502 -3108 2538 -3087
rect 2782 -3108 2818 -3087
rect 2418 -3146 2470 -3136
rect 2418 -3208 2470 -3198
rect 2698 -3146 2750 -3136
rect 2698 -3208 2750 -3198
rect 1730 -3246 1782 -3236
rect 1730 -3308 1782 -3298
rect 2010 -3246 2062 -3236
rect 2010 -3308 2062 -3298
rect 2290 -3246 2342 -3236
rect 2290 -3308 2342 -3298
rect 1662 -3351 1698 -3332
rect 1650 -3357 1708 -3351
rect 1650 -3391 1662 -3357
rect 1696 -3391 1708 -3357
rect 1650 -3397 1708 -3391
rect 1738 -3429 1774 -3308
rect 1942 -3351 1978 -3332
rect 2222 -3351 2258 -3332
rect 1930 -3357 1988 -3351
rect 1930 -3391 1942 -3357
rect 1976 -3391 1988 -3357
rect 1930 -3397 1988 -3391
rect 2210 -3357 2268 -3351
rect 2210 -3391 2222 -3357
rect 2256 -3391 2268 -3357
rect 2210 -3397 2268 -3391
rect 2426 -3429 2462 -3208
rect 2570 -3246 2622 -3236
rect 2570 -3308 2622 -3298
rect 2502 -3351 2538 -3332
rect 2490 -3357 2548 -3351
rect 2490 -3391 2502 -3357
rect 2536 -3391 2548 -3357
rect 2490 -3397 2548 -3391
rect 2578 -3429 2614 -3308
rect 1586 -3441 1658 -3429
rect 1460 -3817 1466 -3490
rect 1420 -3829 1466 -3817
rect 1586 -3817 1618 -3441
rect 1652 -3817 1658 -3441
rect 1586 -3829 1658 -3817
rect 1700 -3441 1774 -3429
rect 1700 -3817 1706 -3441
rect 1740 -3817 1774 -3441
rect 1892 -3441 1938 -3429
rect 1892 -3770 1898 -3441
rect 1700 -3829 1774 -3817
rect 890 -4066 942 -4056
rect 890 -4128 942 -4118
rect 1026 -4156 1062 -3829
rect 1090 -3867 1148 -3861
rect 1090 -3901 1102 -3867
rect 1136 -3901 1148 -3867
rect 1090 -3907 1148 -3901
rect 1102 -3956 1138 -3907
rect 1094 -3966 1146 -3956
rect 1094 -4028 1146 -4018
rect 1178 -4056 1214 -3829
rect 1370 -3867 1428 -3861
rect 1370 -3901 1382 -3867
rect 1416 -3901 1428 -3867
rect 1370 -3907 1428 -3901
rect 1382 -3956 1418 -3907
rect 1374 -3966 1426 -3956
rect 1374 -4028 1426 -4018
rect 1170 -4066 1222 -4056
rect 1170 -4128 1222 -4118
rect 738 -4166 790 -4156
rect 738 -4228 790 -4218
rect 1018 -4166 1070 -4156
rect 1018 -4228 1070 -4218
rect 1178 -4328 1212 -4128
rect 1178 -4358 1418 -4328
rect 1382 -4631 1418 -4358
rect 1586 -4390 1622 -3829
rect 1650 -3867 1708 -3861
rect 1650 -3901 1662 -3867
rect 1696 -3901 1708 -3867
rect 1650 -3907 1708 -3901
rect 1662 -3956 1698 -3907
rect 1654 -3966 1706 -3956
rect 1654 -4028 1706 -4018
rect 1740 -4246 1774 -3829
rect 1866 -3817 1898 -3770
rect 1932 -3817 1938 -3441
rect 1866 -3829 1938 -3817
rect 1980 -3441 2026 -3429
rect 1980 -3817 1986 -3441
rect 2020 -3770 2026 -3441
rect 2172 -3441 2218 -3429
rect 2172 -3770 2178 -3441
rect 2020 -3817 2054 -3770
rect 1980 -3829 2054 -3817
rect 1866 -4156 1902 -3829
rect 1930 -3867 1988 -3861
rect 1930 -3901 1942 -3867
rect 1976 -3901 1988 -3867
rect 1930 -3907 1988 -3901
rect 1942 -3956 1978 -3907
rect 1934 -3966 1986 -3956
rect 1934 -4028 1986 -4018
rect 2018 -4056 2054 -3829
rect 2146 -3817 2178 -3770
rect 2212 -3817 2218 -3441
rect 2146 -3829 2218 -3817
rect 2260 -3441 2306 -3429
rect 2260 -3817 2266 -3441
rect 2300 -3770 2306 -3441
rect 2426 -3441 2498 -3429
rect 2426 -3490 2458 -3441
rect 2300 -3817 2334 -3770
rect 2260 -3829 2334 -3817
rect 2452 -3817 2458 -3490
rect 2492 -3817 2498 -3441
rect 2452 -3829 2498 -3817
rect 2540 -3441 2614 -3429
rect 2540 -3817 2546 -3441
rect 2580 -3490 2614 -3441
rect 2706 -3429 2742 -3208
rect 2850 -3246 2902 -3236
rect 2850 -3308 2902 -3298
rect 2782 -3351 2818 -3332
rect 2770 -3357 2828 -3351
rect 2770 -3391 2782 -3357
rect 2816 -3391 2828 -3357
rect 2770 -3397 2828 -3391
rect 2858 -3429 2894 -3308
rect 2706 -3441 2778 -3429
rect 2706 -3490 2738 -3441
rect 2580 -3817 2586 -3490
rect 2540 -3829 2586 -3817
rect 2732 -3817 2738 -3490
rect 2772 -3817 2778 -3441
rect 2732 -3829 2778 -3817
rect 2820 -3441 2894 -3429
rect 2820 -3817 2826 -3441
rect 2860 -3490 2894 -3441
rect 2860 -3817 2866 -3490
rect 2820 -3829 2866 -3817
rect 2010 -4066 2062 -4056
rect 2010 -4128 2062 -4118
rect 2146 -4156 2182 -3829
rect 2210 -3867 2268 -3861
rect 2210 -3901 2222 -3867
rect 2256 -3901 2268 -3867
rect 2210 -3907 2268 -3901
rect 2222 -3956 2258 -3907
rect 2214 -3966 2266 -3956
rect 2214 -4028 2266 -4018
rect 2298 -4056 2334 -3829
rect 2490 -3867 2548 -3861
rect 2490 -3901 2502 -3867
rect 2536 -3901 2548 -3867
rect 2490 -3907 2548 -3901
rect 2770 -3867 2828 -3861
rect 2770 -3901 2782 -3867
rect 2816 -3901 2828 -3867
rect 2770 -3907 2828 -3901
rect 2502 -3956 2538 -3907
rect 2782 -3956 2818 -3907
rect 2494 -3966 2546 -3956
rect 2494 -4028 2546 -4018
rect 2774 -3966 2826 -3956
rect 2774 -4028 2826 -4018
rect 2290 -4066 2342 -4056
rect 2290 -4128 2342 -4118
rect 1858 -4166 1910 -4156
rect 1858 -4228 1910 -4218
rect 2138 -4166 2190 -4156
rect 2138 -4228 2190 -4218
rect 1458 -4426 1622 -4390
rect 1662 -4276 1774 -4246
rect 1458 -4428 1510 -4426
rect 1458 -4490 1510 -4480
rect 1370 -4637 1428 -4631
rect 1370 -4671 1382 -4637
rect 1416 -4671 1428 -4637
rect 1370 -4677 1428 -4671
rect 1458 -4709 1494 -4490
rect 1578 -4520 1630 -4510
rect 1578 -4582 1630 -4572
rect 1332 -4721 1378 -4709
rect 1332 -5068 1338 -4721
rect 1304 -5097 1338 -5068
rect 1372 -5097 1378 -4721
rect 1304 -5109 1378 -5097
rect 1420 -4721 1494 -4709
rect 1420 -5097 1426 -4721
rect 1460 -4802 1494 -4721
rect 1584 -4709 1620 -4582
rect 1662 -4631 1698 -4276
rect 2148 -4338 2182 -4228
rect 1740 -4376 2182 -4338
rect 1650 -4637 1708 -4631
rect 1650 -4671 1662 -4637
rect 1696 -4671 1708 -4637
rect 1650 -4677 1708 -4671
rect 1740 -4709 1776 -4376
rect 1584 -4721 1658 -4709
rect 1460 -5097 1466 -4802
rect 1584 -4804 1618 -4721
rect 1420 -5109 1466 -5097
rect 1612 -5097 1618 -4804
rect 1652 -5097 1658 -4721
rect 1612 -5109 1658 -5097
rect 1700 -4721 1776 -4709
rect 1700 -5097 1706 -4721
rect 1740 -5097 1776 -4721
rect 1700 -5109 1776 -5097
rect 1304 -5338 1340 -5109
rect 1370 -5147 1428 -5141
rect 1370 -5181 1382 -5147
rect 1416 -5181 1428 -5147
rect 1650 -5147 1708 -5141
rect 1650 -5148 1662 -5147
rect 1370 -5187 1428 -5181
rect 1480 -5181 1662 -5148
rect 1696 -5181 1708 -5147
rect 1480 -5182 1708 -5181
rect 1382 -5234 1418 -5187
rect 1374 -5244 1426 -5234
rect 1374 -5306 1426 -5296
rect 1296 -5348 1348 -5338
rect 1480 -5342 1514 -5182
rect 1650 -5187 1708 -5182
rect 1654 -5244 1706 -5234
rect 1654 -5306 1706 -5296
rect 1296 -5410 1348 -5400
rect 1382 -5376 1514 -5342
rect 1382 -5489 1418 -5376
rect 1458 -5428 1510 -5418
rect 1369 -5495 1427 -5489
rect 1369 -5529 1381 -5495
rect 1415 -5529 1427 -5495
rect 1369 -5535 1427 -5529
rect 1458 -5490 1510 -5480
rect 1662 -5489 1698 -5306
rect 1740 -5324 1776 -5109
rect 1804 -4428 1856 -4418
rect 1804 -4486 1856 -4480
rect 1804 -5296 1854 -4486
rect 1734 -5334 1786 -5324
rect 1734 -5396 1786 -5386
rect 1814 -5424 1854 -5296
rect 1458 -5567 1494 -5490
rect 1649 -5495 1707 -5489
rect 1649 -5529 1661 -5495
rect 1695 -5529 1707 -5495
rect 1649 -5535 1707 -5529
rect 1331 -5579 1377 -5567
rect 1331 -5955 1337 -5579
rect 1371 -5955 1377 -5579
rect 1331 -5967 1377 -5955
rect 1419 -5579 1494 -5567
rect 1419 -5955 1425 -5579
rect 1459 -5606 1494 -5579
rect 1611 -5579 1657 -5567
rect 1459 -5955 1465 -5606
rect 1611 -5792 1617 -5579
rect 1419 -5967 1465 -5955
rect 1584 -5955 1617 -5792
rect 1651 -5955 1657 -5579
rect 1584 -5967 1657 -5955
rect 1699 -5579 1745 -5567
rect 1699 -5955 1705 -5579
rect 1739 -5955 1745 -5579
rect 1699 -5967 1745 -5955
rect 154 -6156 254 -6056
rect 1338 -6124 1374 -5967
rect 1584 -6028 1620 -5967
rect 1706 -6004 1742 -5967
rect 1804 -6004 1854 -5424
rect 1576 -6038 1628 -6028
rect 1706 -6040 1854 -6004
rect 1576 -6100 1628 -6090
rect 1330 -6134 1382 -6124
rect 190 -6224 218 -6156
rect 1584 -6150 1620 -6100
rect 2576 -6134 2628 -6124
rect 1584 -6182 2342 -6150
rect 1330 -6196 1382 -6186
rect 150 -6252 2114 -6224
rect 150 -8016 178 -6252
rect 254 -6324 306 -6314
rect 254 -6386 306 -6376
rect 534 -6324 586 -6314
rect 534 -6386 586 -6376
rect 262 -6434 298 -6386
rect 542 -6434 578 -6386
rect 250 -6440 308 -6434
rect 250 -6474 262 -6440
rect 296 -6474 308 -6440
rect 250 -6480 308 -6474
rect 530 -6440 588 -6434
rect 530 -6474 542 -6440
rect 576 -6474 588 -6440
rect 530 -6480 588 -6474
rect 810 -6440 868 -6434
rect 966 -6440 994 -6252
rect 1374 -6324 1426 -6314
rect 1374 -6386 1426 -6376
rect 1654 -6324 1706 -6314
rect 1654 -6386 1706 -6376
rect 1382 -6434 1418 -6386
rect 1662 -6434 1698 -6386
rect 1090 -6440 1148 -6434
rect 810 -6474 822 -6440
rect 856 -6474 1102 -6440
rect 1136 -6474 1148 -6440
rect 810 -6476 1148 -6474
rect 810 -6480 868 -6476
rect 1090 -6480 1148 -6476
rect 1370 -6440 1428 -6434
rect 1370 -6474 1382 -6440
rect 1416 -6474 1428 -6440
rect 1370 -6480 1428 -6474
rect 1650 -6440 1708 -6434
rect 1650 -6474 1662 -6440
rect 1696 -6474 1708 -6440
rect 1650 -6480 1708 -6474
rect 1930 -6440 1988 -6434
rect 2086 -6440 2114 -6252
rect 2210 -6440 2268 -6434
rect 1930 -6474 1942 -6440
rect 1976 -6474 2222 -6440
rect 2256 -6474 2268 -6440
rect 1930 -6476 2268 -6474
rect 1930 -6480 1988 -6476
rect 2210 -6480 2268 -6476
rect 2306 -6512 2342 -6182
rect 2576 -6196 2628 -6186
rect 2494 -6324 2546 -6314
rect 2494 -6386 2546 -6376
rect 2502 -6434 2538 -6386
rect 2490 -6440 2548 -6434
rect 2490 -6474 2502 -6440
rect 2536 -6474 2548 -6440
rect 2490 -6480 2548 -6474
rect 2586 -6512 2624 -6196
rect 2750 -6256 2850 -6156
rect 2782 -6314 2816 -6256
rect 2774 -6324 2826 -6314
rect 2774 -6386 2826 -6376
rect 2782 -6434 2818 -6386
rect 2770 -6440 2828 -6434
rect 2770 -6474 2782 -6440
rect 2816 -6474 2828 -6440
rect 2770 -6480 2828 -6474
rect 212 -6524 258 -6512
rect 212 -6900 218 -6524
rect 252 -6900 258 -6524
rect 212 -6912 258 -6900
rect 300 -6524 346 -6512
rect 300 -6900 306 -6524
rect 340 -6682 346 -6524
rect 492 -6524 538 -6512
rect 340 -6900 382 -6682
rect 300 -6912 382 -6900
rect 212 -7020 246 -6912
rect 346 -6948 382 -6912
rect 492 -6900 498 -6524
rect 532 -6900 538 -6524
rect 492 -6912 538 -6900
rect 580 -6524 626 -6512
rect 580 -6900 586 -6524
rect 620 -6682 626 -6524
rect 772 -6524 818 -6512
rect 620 -6900 662 -6682
rect 580 -6912 662 -6900
rect 338 -6958 390 -6948
rect 338 -7020 390 -7010
rect 212 -7030 298 -7020
rect 212 -7082 246 -7030
rect 212 -7092 298 -7082
rect 492 -7028 526 -6912
rect 626 -6948 662 -6912
rect 772 -6900 778 -6524
rect 812 -6900 818 -6524
rect 772 -6912 818 -6900
rect 860 -6524 906 -6512
rect 860 -6900 866 -6524
rect 900 -6682 906 -6524
rect 1052 -6524 1098 -6512
rect 900 -6900 942 -6682
rect 860 -6912 942 -6900
rect 618 -6958 670 -6948
rect 618 -7020 670 -7010
rect 772 -7028 806 -6912
rect 492 -7038 544 -7028
rect 212 -7210 246 -7092
rect 492 -7100 544 -7090
rect 772 -7038 824 -7028
rect 772 -7100 824 -7090
rect 338 -7114 390 -7104
rect 338 -7176 390 -7166
rect 346 -7210 382 -7176
rect 212 -7222 258 -7210
rect 212 -7598 218 -7222
rect 252 -7598 258 -7222
rect 212 -7610 258 -7598
rect 300 -7222 382 -7210
rect 300 -7598 306 -7222
rect 340 -7442 382 -7222
rect 492 -7210 526 -7100
rect 618 -7114 670 -7104
rect 618 -7176 670 -7166
rect 626 -7210 662 -7176
rect 492 -7222 538 -7210
rect 340 -7598 346 -7442
rect 300 -7610 346 -7598
rect 492 -7598 498 -7222
rect 532 -7598 538 -7222
rect 492 -7610 538 -7598
rect 580 -7222 662 -7210
rect 580 -7598 586 -7222
rect 620 -7442 662 -7222
rect 772 -7210 806 -7100
rect 906 -7104 942 -6912
rect 1052 -6900 1058 -6524
rect 1092 -6900 1098 -6524
rect 1052 -6912 1098 -6900
rect 1140 -6524 1186 -6512
rect 1140 -6900 1146 -6524
rect 1180 -6682 1186 -6524
rect 1332 -6524 1378 -6512
rect 1180 -6900 1222 -6682
rect 1140 -6912 1222 -6900
rect 1052 -7028 1086 -6912
rect 1052 -7038 1104 -7028
rect 1052 -7100 1104 -7090
rect 898 -7114 950 -7104
rect 898 -7176 950 -7166
rect 1052 -7210 1086 -7100
rect 1186 -7104 1222 -6912
rect 1332 -6900 1338 -6524
rect 1372 -6900 1378 -6524
rect 1332 -6912 1378 -6900
rect 1420 -6524 1466 -6512
rect 1420 -6900 1426 -6524
rect 1460 -6682 1466 -6524
rect 1612 -6524 1658 -6512
rect 1460 -6900 1502 -6682
rect 1420 -6912 1502 -6900
rect 1332 -7028 1366 -6912
rect 1466 -6948 1502 -6912
rect 1612 -6900 1618 -6524
rect 1652 -6900 1658 -6524
rect 1612 -6912 1658 -6900
rect 1700 -6524 1746 -6512
rect 1700 -6900 1706 -6524
rect 1740 -6682 1746 -6524
rect 1892 -6524 1938 -6512
rect 1740 -6900 1782 -6682
rect 1700 -6912 1782 -6900
rect 1458 -6958 1510 -6948
rect 1458 -7020 1510 -7010
rect 1612 -7028 1646 -6912
rect 1746 -6948 1782 -6912
rect 1892 -6900 1898 -6524
rect 1932 -6900 1938 -6524
rect 1892 -6912 1938 -6900
rect 1980 -6524 2026 -6512
rect 1980 -6900 1986 -6524
rect 2020 -6682 2026 -6524
rect 2172 -6524 2218 -6512
rect 2020 -6900 2062 -6682
rect 1980 -6912 2062 -6900
rect 1738 -6958 1790 -6948
rect 1738 -7020 1790 -7010
rect 1892 -7028 1926 -6912
rect 1332 -7038 1384 -7028
rect 1332 -7100 1384 -7090
rect 1612 -7038 1664 -7028
rect 1612 -7100 1664 -7090
rect 1892 -7038 1944 -7028
rect 1892 -7100 1944 -7090
rect 1178 -7114 1230 -7104
rect 1178 -7176 1230 -7166
rect 1332 -7210 1366 -7100
rect 1458 -7114 1510 -7104
rect 1458 -7176 1510 -7166
rect 1466 -7210 1502 -7176
rect 772 -7222 818 -7210
rect 620 -7598 626 -7442
rect 580 -7610 626 -7598
rect 772 -7598 778 -7222
rect 812 -7598 818 -7222
rect 772 -7610 818 -7598
rect 860 -7222 906 -7210
rect 860 -7598 866 -7222
rect 900 -7442 906 -7222
rect 1052 -7222 1098 -7210
rect 900 -7598 942 -7442
rect 860 -7610 942 -7598
rect 1052 -7598 1058 -7222
rect 1092 -7598 1098 -7222
rect 1052 -7610 1098 -7598
rect 1140 -7222 1186 -7210
rect 1140 -7598 1146 -7222
rect 1180 -7442 1186 -7222
rect 1332 -7222 1378 -7210
rect 1180 -7598 1222 -7442
rect 1140 -7610 1222 -7598
rect 1332 -7598 1338 -7222
rect 1372 -7598 1378 -7222
rect 1332 -7610 1378 -7598
rect 1420 -7222 1502 -7210
rect 1420 -7598 1426 -7222
rect 1460 -7442 1502 -7222
rect 1612 -7210 1646 -7100
rect 1738 -7114 1790 -7104
rect 1738 -7176 1790 -7166
rect 1746 -7210 1782 -7176
rect 1612 -7222 1658 -7210
rect 1460 -7598 1466 -7442
rect 1420 -7610 1466 -7598
rect 1612 -7598 1618 -7222
rect 1652 -7598 1658 -7222
rect 1612 -7610 1658 -7598
rect 1700 -7222 1782 -7210
rect 1700 -7598 1706 -7222
rect 1740 -7442 1782 -7222
rect 1892 -7210 1926 -7100
rect 2026 -7104 2062 -6912
rect 2172 -6900 2178 -6524
rect 2212 -6900 2218 -6524
rect 2172 -6912 2218 -6900
rect 2260 -6524 2342 -6512
rect 2260 -6900 2266 -6524
rect 2300 -6900 2342 -6524
rect 2260 -6912 2342 -6900
rect 2172 -7028 2206 -6912
rect 2172 -7038 2224 -7028
rect 2172 -7100 2224 -7090
rect 2018 -7114 2070 -7104
rect 2018 -7176 2070 -7166
rect 2172 -7210 2206 -7100
rect 2306 -7104 2342 -6912
rect 2452 -6524 2498 -6512
rect 2452 -6900 2458 -6524
rect 2492 -6900 2498 -6524
rect 2452 -6912 2498 -6900
rect 2540 -6524 2624 -6512
rect 2540 -6900 2546 -6524
rect 2580 -6732 2624 -6524
rect 2732 -6524 2778 -6512
rect 2580 -6900 2622 -6732
rect 2540 -6912 2622 -6900
rect 2452 -7028 2486 -6912
rect 2586 -6948 2622 -6912
rect 2732 -6900 2738 -6524
rect 2772 -6900 2778 -6524
rect 2732 -6912 2778 -6900
rect 2820 -6524 2866 -6512
rect 2820 -6900 2826 -6524
rect 2860 -6682 2866 -6524
rect 2860 -6900 2902 -6682
rect 2820 -6912 2902 -6900
rect 2578 -6958 2630 -6948
rect 2578 -7020 2630 -7010
rect 2452 -7038 2504 -7028
rect 2732 -7048 2766 -6912
rect 2866 -6948 2902 -6912
rect 2858 -6958 2910 -6948
rect 2858 -7020 2910 -7010
rect 3184 -7048 3284 -7020
rect 3628 -7048 3634 -2410
rect 2504 -7076 3634 -7048
rect 2452 -7100 2504 -7090
rect 2298 -7114 2350 -7104
rect 2298 -7176 2350 -7166
rect 2452 -7210 2486 -7100
rect 2578 -7114 2630 -7104
rect 2578 -7176 2630 -7166
rect 2586 -7210 2622 -7176
rect 1892 -7222 1938 -7210
rect 1740 -7598 1746 -7442
rect 1700 -7610 1746 -7598
rect 1892 -7598 1898 -7222
rect 1932 -7598 1938 -7222
rect 1892 -7610 1938 -7598
rect 1980 -7222 2026 -7210
rect 1980 -7598 1986 -7222
rect 2020 -7442 2026 -7222
rect 2172 -7222 2218 -7210
rect 2020 -7598 2062 -7442
rect 1980 -7610 2062 -7598
rect 2172 -7598 2178 -7222
rect 2212 -7598 2218 -7222
rect 2172 -7610 2218 -7598
rect 2260 -7222 2306 -7210
rect 2260 -7598 2266 -7222
rect 2300 -7442 2306 -7222
rect 2452 -7222 2498 -7210
rect 2300 -7598 2342 -7442
rect 2260 -7610 2342 -7598
rect 2452 -7598 2458 -7222
rect 2492 -7598 2498 -7222
rect 2452 -7610 2498 -7598
rect 2540 -7222 2622 -7210
rect 2540 -7598 2546 -7222
rect 2580 -7442 2622 -7222
rect 2732 -7210 2766 -7076
rect 2858 -7114 2910 -7104
rect 3184 -7120 3284 -7076
rect 2858 -7176 2910 -7166
rect 2866 -7210 2902 -7176
rect 2732 -7222 2778 -7210
rect 2580 -7598 2586 -7442
rect 2540 -7610 2586 -7598
rect 2732 -7598 2738 -7222
rect 2772 -7598 2778 -7222
rect 2732 -7610 2778 -7598
rect 2820 -7222 2902 -7210
rect 2820 -7598 2826 -7222
rect 2860 -7442 2902 -7222
rect 2860 -7598 2866 -7442
rect 2820 -7610 2866 -7598
rect 250 -7648 588 -7642
rect 250 -7682 262 -7648
rect 296 -7682 542 -7648
rect 576 -7682 588 -7648
rect 250 -7688 588 -7682
rect 810 -7648 868 -7642
rect 810 -7682 822 -7648
rect 856 -7682 868 -7648
rect 810 -7688 868 -7682
rect 406 -8016 434 -7688
rect 822 -7738 858 -7688
rect 814 -7748 866 -7738
rect 814 -7810 866 -7800
rect 906 -7832 942 -7610
rect 1090 -7648 1148 -7642
rect 1090 -7682 1102 -7648
rect 1136 -7682 1148 -7648
rect 1090 -7688 1148 -7682
rect 1102 -7738 1138 -7688
rect 1094 -7748 1146 -7738
rect 1094 -7810 1146 -7800
rect 1186 -7832 1222 -7610
rect 1370 -7648 1428 -7642
rect 1650 -7648 1708 -7642
rect 1370 -7682 1382 -7648
rect 1416 -7682 1662 -7648
rect 1696 -7682 1708 -7648
rect 1370 -7684 1708 -7682
rect 1370 -7688 1428 -7684
rect 898 -7842 950 -7832
rect 898 -7904 950 -7894
rect 1178 -7842 1230 -7832
rect 1178 -7904 1230 -7894
rect 1526 -8016 1554 -7684
rect 1650 -7688 1708 -7684
rect 1930 -7648 1988 -7642
rect 1930 -7682 1942 -7648
rect 1976 -7682 1988 -7648
rect 1930 -7688 1988 -7682
rect 1934 -7748 1986 -7688
rect 1934 -7810 1986 -7800
rect 2026 -7832 2062 -7610
rect 2210 -7648 2268 -7642
rect 2210 -7682 2222 -7648
rect 2256 -7682 2268 -7648
rect 2210 -7688 2268 -7682
rect 2222 -7738 2258 -7688
rect 2214 -7748 2266 -7738
rect 2214 -7810 2266 -7800
rect 2306 -7832 2342 -7610
rect 2490 -7648 2548 -7642
rect 2770 -7648 2828 -7642
rect 2490 -7682 2502 -7648
rect 2536 -7682 2782 -7648
rect 2816 -7682 2828 -7648
rect 2490 -7684 2828 -7682
rect 2490 -7688 2548 -7684
rect 2018 -7842 2070 -7832
rect 2018 -7904 2070 -7894
rect 2298 -7842 2350 -7832
rect 2298 -7904 2350 -7894
rect 2646 -8016 2674 -7684
rect 2770 -7688 2828 -7684
rect 150 -8044 2674 -8016
rect -502 -8488 -390 -8162
rect 3628 -8162 3634 -7076
rect 3734 -8162 3740 -2410
rect 210 -8488 220 -8188
rect 3018 -8488 3028 -8188
rect 3628 -8488 3740 -8162
rect -502 -8494 3740 -8488
rect -502 -8594 -396 -8494
rect 3634 -8594 3740 -8494
rect -502 -8600 3740 -8594
<< via1 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -110 440 -58 492
rect 170 440 222 492
rect -26 346 26 398
rect 450 440 502 492
rect 254 346 306 398
rect 730 440 782 492
rect 534 346 586 398
rect 1010 440 1062 492
rect 814 346 866 398
rect 1290 440 1342 492
rect 1094 346 1146 398
rect 1570 440 1622 492
rect 1374 346 1426 398
rect 1850 440 1902 492
rect 1654 346 1706 398
rect 2130 440 2182 492
rect 1934 346 1986 398
rect 2410 440 2462 492
rect 2214 346 2266 398
rect 2690 440 2742 492
rect 2494 346 2546 398
rect 2970 440 3022 492
rect 2774 346 2826 398
rect 3238 238 3290 290
rect 60 -382 112 -330
rect 340 -382 392 -330
rect 620 -382 672 -330
rect 900 -382 952 -330
rect 1180 -382 1232 -330
rect 1460 -382 1512 -330
rect 1740 -382 1792 -330
rect 2020 -382 2072 -330
rect 2300 -382 2352 -330
rect 2580 -382 2632 -330
rect 2860 -382 2912 -330
rect 3140 -382 3192 -330
rect -26 -1114 26 -1062
rect 254 -1114 306 -1062
rect 534 -1114 586 -1062
rect 814 -1114 866 -1062
rect 1094 -1114 1146 -1062
rect 1934 -1114 1986 -1062
rect 2214 -1114 2266 -1062
rect 2494 -1114 2546 -1062
rect 2774 -1114 2826 -1062
rect 3054 -1114 3106 -1062
rect 1374 -1230 1426 -1178
rect 1654 -1230 1706 -1178
rect 414 -1514 466 -1462
rect 2478 -1424 2530 -1372
rect 2916 -1862 2968 -1810
rect 900 -2194 952 -2142
rect 2774 -2186 2826 -2134
rect 330 -2274 382 -2222
rect 610 -2274 662 -2222
rect 178 -2374 230 -2322
rect 254 -2474 306 -2422
rect 458 -2374 510 -2322
rect 534 -2474 586 -2422
rect 814 -2474 866 -2422
rect 1450 -2274 1502 -2222
rect 1730 -2274 1782 -2222
rect 2570 -2274 2622 -2222
rect 1298 -2374 1350 -2322
rect 1094 -2474 1146 -2422
rect 1374 -2474 1426 -2422
rect 1578 -2374 1630 -2322
rect 1654 -2474 1706 -2422
rect 2418 -2374 2470 -2322
rect 1934 -2474 1986 -2422
rect 2214 -2474 2266 -2422
rect 2494 -2474 2546 -2422
rect 2698 -2374 2750 -2322
rect 178 -3198 230 -3146
rect 458 -3198 510 -3146
rect 738 -3194 790 -3142
rect 330 -3298 382 -3246
rect 1018 -3194 1070 -3142
rect 1298 -3198 1350 -3146
rect 1578 -3198 1630 -3146
rect 1858 -3194 1910 -3142
rect 610 -3298 662 -3246
rect 890 -3298 942 -3246
rect 1170 -3298 1222 -3246
rect 1450 -3298 1502 -3246
rect 254 -4018 306 -3966
rect 534 -4018 586 -3966
rect 814 -4018 866 -3966
rect 2850 -2274 2902 -2222
rect 2774 -2474 2826 -2422
rect 2138 -3194 2190 -3142
rect 2418 -3198 2470 -3146
rect 2698 -3198 2750 -3146
rect 1730 -3298 1782 -3246
rect 2010 -3298 2062 -3246
rect 2290 -3298 2342 -3246
rect 2570 -3298 2622 -3246
rect 890 -4118 942 -4066
rect 1094 -4018 1146 -3966
rect 1374 -4018 1426 -3966
rect 1170 -4118 1222 -4066
rect 738 -4218 790 -4166
rect 1018 -4218 1070 -4166
rect 1654 -4018 1706 -3966
rect 1934 -4018 1986 -3966
rect 2850 -3298 2902 -3246
rect 2010 -4118 2062 -4066
rect 2214 -4018 2266 -3966
rect 2494 -4018 2546 -3966
rect 2774 -4018 2826 -3966
rect 2290 -4118 2342 -4066
rect 1858 -4218 1910 -4166
rect 2138 -4218 2190 -4166
rect 1458 -4480 1510 -4428
rect 1578 -4572 1630 -4520
rect 1374 -5296 1426 -5244
rect 1654 -5296 1706 -5244
rect 1296 -5400 1348 -5348
rect 1458 -5480 1510 -5428
rect 1804 -4480 1856 -4428
rect 1734 -5386 1786 -5334
rect 1576 -6090 1628 -6038
rect 1330 -6186 1382 -6134
rect 254 -6376 306 -6324
rect 534 -6376 586 -6324
rect 1374 -6376 1426 -6324
rect 1654 -6376 1706 -6324
rect 2576 -6186 2628 -6134
rect 2494 -6376 2546 -6324
rect 2774 -6376 2826 -6324
rect 338 -7010 390 -6958
rect 246 -7082 298 -7030
rect 618 -7010 670 -6958
rect 492 -7090 544 -7038
rect 772 -7090 824 -7038
rect 338 -7166 390 -7114
rect 618 -7166 670 -7114
rect 1052 -7090 1104 -7038
rect 898 -7166 950 -7114
rect 1458 -7010 1510 -6958
rect 1738 -7010 1790 -6958
rect 1332 -7090 1384 -7038
rect 1612 -7090 1664 -7038
rect 1892 -7090 1944 -7038
rect 1178 -7166 1230 -7114
rect 1458 -7166 1510 -7114
rect 1738 -7166 1790 -7114
rect 2172 -7090 2224 -7038
rect 2018 -7166 2070 -7114
rect 2578 -7010 2630 -6958
rect 2452 -7090 2504 -7038
rect 2858 -7010 2910 -6958
rect 2298 -7166 2350 -7114
rect 2578 -7166 2630 -7114
rect 2858 -7166 2910 -7114
rect 814 -7800 866 -7748
rect 1094 -7800 1146 -7748
rect 898 -7894 950 -7842
rect 1178 -7894 1230 -7842
rect 1934 -7800 1986 -7748
rect 2214 -7800 2266 -7748
rect 2018 -7894 2070 -7842
rect 2298 -7894 2350 -7842
rect -390 -8488 210 -8188
rect 3028 -8488 3628 -8188
<< metal2 >>
rect -390 1016 210 1026
rect -390 706 210 716
rect 3028 1016 3628 1026
rect 3028 706 3628 716
rect -120 440 -110 492
rect -58 440 170 492
rect 222 440 450 492
rect 502 440 730 492
rect 782 440 1010 492
rect 1062 440 1290 492
rect 1342 440 1570 492
rect 1622 440 1850 492
rect 1902 440 2130 492
rect 2182 440 2410 492
rect 2462 440 2690 492
rect 2742 440 2970 492
rect 3022 440 3032 492
rect -190 346 -26 398
rect 26 346 36 398
rect 244 346 254 398
rect 306 396 316 398
rect 524 396 534 398
rect 306 346 534 396
rect 586 396 596 398
rect 804 396 814 398
rect 586 346 814 396
rect 866 396 876 398
rect 1084 396 1094 398
rect 866 346 1094 396
rect 1146 396 1156 398
rect 1364 396 1374 398
rect 1146 346 1374 396
rect 1426 396 1436 398
rect 1644 396 1654 398
rect 1426 346 1654 396
rect 1706 396 1716 398
rect 1924 396 1934 398
rect 1706 346 1934 396
rect 1986 396 1996 398
rect 2204 396 2214 398
rect 1986 346 2214 396
rect 2266 396 2276 398
rect 2484 396 2494 398
rect 2266 346 2494 396
rect 2546 396 2556 398
rect 2764 396 2774 398
rect 2546 346 2774 396
rect 2826 396 2836 398
rect 3338 396 3390 398
rect 2826 346 3390 396
rect -190 -1178 -138 346
rect 3238 290 3290 300
rect 50 -382 60 -330
rect 112 -382 340 -330
rect 392 -382 620 -330
rect 672 -382 900 -330
rect 952 -382 1180 -330
rect 1232 -382 1460 -330
rect 1512 -382 1522 -330
rect 1730 -382 1740 -330
rect 1792 -382 2020 -330
rect 2072 -382 2300 -330
rect 2352 -382 2580 -330
rect 2632 -382 2860 -330
rect 2912 -382 3140 -330
rect 3192 -382 3202 -330
rect -36 -1114 -26 -1062
rect 26 -1114 254 -1062
rect 306 -1114 534 -1062
rect 586 -1114 814 -1062
rect 866 -1114 1094 -1062
rect 1146 -1114 1934 -1062
rect 1986 -1114 2214 -1062
rect 2266 -1114 2494 -1062
rect 2546 -1114 2774 -1062
rect 2826 -1114 3054 -1062
rect 3106 -1114 3116 -1062
rect -190 -1230 1374 -1178
rect 1426 -1230 1436 -1178
rect 414 -1462 466 -1452
rect 414 -1764 466 -1514
rect 964 -1466 1016 -1230
rect 1514 -1258 1566 -1114
rect 3238 -1178 3290 238
rect 1644 -1230 1654 -1178
rect 1706 -1230 3290 -1178
rect 3338 -1258 3390 346
rect 1514 -1310 3390 -1258
rect 2478 -1372 2530 -1362
rect 1954 -1466 2000 -1464
rect 2478 -1466 2530 -1424
rect 964 -1518 2530 -1466
rect 414 -1804 806 -1764
rect 774 -2154 806 -1804
rect 890 -2154 900 -2142
rect 774 -2194 900 -2154
rect 952 -2194 962 -2142
rect 1954 -2222 2000 -1518
rect 2916 -1810 2972 -1310
rect 2968 -1862 2972 -1810
rect 2916 -2134 2972 -1862
rect 2764 -2186 2774 -2134
rect 2826 -2186 2972 -2134
rect 2916 -2188 2972 -2186
rect 320 -2274 330 -2222
rect 382 -2274 610 -2222
rect 662 -2274 1450 -2222
rect 1502 -2274 1730 -2222
rect 1782 -2274 2570 -2222
rect 2622 -2274 2850 -2222
rect 2902 -2274 3104 -2222
rect -76 -2374 178 -2322
rect 230 -2374 458 -2322
rect 510 -2374 1298 -2322
rect 1350 -2374 1578 -2322
rect 1630 -2374 2418 -2322
rect 2470 -2374 2698 -2322
rect 2750 -2374 2760 -2322
rect -76 -4166 -24 -2374
rect 58 -2474 254 -2422
rect 306 -2474 534 -2422
rect 586 -2474 814 -2422
rect 866 -2474 1094 -2422
rect 1146 -2474 1374 -2422
rect 1426 -2474 1654 -2422
rect 1706 -2474 1934 -2422
rect 1986 -2474 2214 -2422
rect 2266 -2474 2494 -2422
rect 2546 -2474 2774 -2422
rect 2826 -2474 3022 -2422
rect 58 -3966 110 -2474
rect 728 -3146 738 -3142
rect 168 -3198 178 -3146
rect 230 -3198 458 -3146
rect 510 -3194 738 -3146
rect 790 -3146 800 -3142
rect 1008 -3146 1018 -3142
rect 790 -3194 1018 -3146
rect 1070 -3146 1080 -3142
rect 1848 -3146 1858 -3142
rect 1070 -3194 1298 -3146
rect 510 -3198 1298 -3194
rect 1350 -3198 1578 -3146
rect 1630 -3194 1858 -3146
rect 1910 -3146 1920 -3142
rect 2128 -3146 2138 -3142
rect 1910 -3194 2138 -3146
rect 2190 -3146 2200 -3142
rect 2190 -3194 2418 -3146
rect 1630 -3198 2418 -3194
rect 2470 -3198 2698 -3146
rect 2750 -3198 2760 -3146
rect 320 -3298 330 -3246
rect 382 -3298 610 -3246
rect 662 -3298 890 -3246
rect 942 -3298 1170 -3246
rect 1222 -3298 1450 -3246
rect 1502 -3298 1730 -3246
rect 1782 -3298 2010 -3246
rect 2062 -3298 2290 -3246
rect 2342 -3298 2570 -3246
rect 2622 -3298 2850 -3246
rect 2902 -3298 2912 -3246
rect 330 -3300 2902 -3298
rect 2970 -3966 3022 -2474
rect 58 -4018 254 -3966
rect 306 -4018 534 -3966
rect 586 -4018 814 -3966
rect 866 -4018 1094 -3966
rect 1146 -4018 1374 -3966
rect 1426 -4018 1654 -3966
rect 1706 -4018 1934 -3966
rect 1986 -4018 2214 -3966
rect 2266 -4018 2494 -3966
rect 2546 -4018 2774 -3966
rect 2826 -4018 3022 -3966
rect 3052 -4066 3104 -2274
rect 880 -4118 890 -4066
rect 942 -4118 1170 -4066
rect 1222 -4118 2010 -4066
rect 2062 -4118 2290 -4066
rect 2342 -4118 3104 -4066
rect -76 -4218 738 -4166
rect 790 -4218 1018 -4166
rect 1070 -4218 1858 -4166
rect 1910 -4218 2138 -4166
rect 2190 -4218 2200 -4166
rect 1448 -4480 1458 -4428
rect 1510 -4480 1804 -4428
rect 1856 -4480 1866 -4428
rect 1568 -4572 1578 -4520
rect 1630 -4572 1876 -4520
rect 1364 -5296 1374 -5244
rect 1426 -5296 1654 -5244
rect 1706 -5296 1716 -5244
rect 1724 -5346 1734 -5334
rect 1286 -5400 1296 -5348
rect 1348 -5400 1358 -5348
rect 1554 -5380 1734 -5346
rect 1296 -6038 1348 -5400
rect 1554 -5428 1588 -5380
rect 1724 -5386 1734 -5380
rect 1786 -5386 1796 -5334
rect 1448 -5480 1458 -5428
rect 1510 -5480 1588 -5428
rect 1296 -6090 1576 -6038
rect 1628 -6090 1638 -6038
rect 1826 -6134 1876 -4572
rect 1320 -6186 1330 -6134
rect 1382 -6186 2576 -6134
rect 2628 -6186 2638 -6134
rect 138 -6376 254 -6324
rect 306 -6376 534 -6324
rect 586 -6376 1374 -6324
rect 1426 -6376 1654 -6324
rect 1706 -6376 2494 -6324
rect 2546 -6376 2774 -6324
rect 2826 -6376 2836 -6324
rect 138 -7748 196 -6376
rect 328 -7010 338 -6958
rect 390 -7010 618 -6958
rect 670 -7010 1458 -6958
rect 1510 -7010 1738 -6958
rect 1790 -7010 2578 -6958
rect 2630 -7010 2858 -6958
rect 2910 -7010 3026 -6958
rect 236 -7082 246 -7030
rect 298 -7048 308 -7030
rect 482 -7048 492 -7038
rect 298 -7076 492 -7048
rect 298 -7082 308 -7076
rect 482 -7090 492 -7076
rect 544 -7048 554 -7038
rect 762 -7048 772 -7038
rect 544 -7076 772 -7048
rect 544 -7090 554 -7076
rect 762 -7090 772 -7076
rect 824 -7048 834 -7038
rect 1042 -7048 1052 -7038
rect 824 -7076 1052 -7048
rect 824 -7090 834 -7076
rect 1042 -7090 1052 -7076
rect 1104 -7048 1114 -7038
rect 1322 -7048 1332 -7038
rect 1104 -7076 1332 -7048
rect 1104 -7090 1114 -7076
rect 1322 -7090 1332 -7076
rect 1384 -7048 1394 -7038
rect 1602 -7048 1612 -7038
rect 1384 -7076 1612 -7048
rect 1384 -7090 1394 -7076
rect 1602 -7090 1612 -7076
rect 1664 -7048 1674 -7038
rect 1882 -7048 1892 -7038
rect 1664 -7076 1892 -7048
rect 1664 -7090 1674 -7076
rect 1882 -7090 1892 -7076
rect 1944 -7048 1954 -7038
rect 2162 -7048 2172 -7038
rect 1944 -7076 2172 -7048
rect 1944 -7090 1954 -7076
rect 2162 -7090 2172 -7076
rect 2224 -7048 2234 -7038
rect 2442 -7048 2452 -7038
rect 2224 -7076 2452 -7048
rect 2224 -7090 2234 -7076
rect 2442 -7090 2452 -7076
rect 2504 -7090 2514 -7038
rect 328 -7166 338 -7114
rect 390 -7118 396 -7114
rect 612 -7118 618 -7114
rect 390 -7166 618 -7118
rect 670 -7118 676 -7114
rect 892 -7118 898 -7114
rect 670 -7166 898 -7118
rect 950 -7118 956 -7114
rect 1172 -7118 1178 -7114
rect 950 -7166 1178 -7118
rect 1230 -7118 1236 -7114
rect 1452 -7118 1458 -7114
rect 1230 -7166 1458 -7118
rect 1510 -7118 1516 -7114
rect 1732 -7118 1738 -7114
rect 1510 -7166 1738 -7118
rect 1790 -7118 1796 -7114
rect 2012 -7118 2018 -7114
rect 1790 -7166 2018 -7118
rect 2070 -7118 2076 -7114
rect 2292 -7118 2298 -7114
rect 2070 -7166 2298 -7118
rect 2350 -7118 2356 -7114
rect 2572 -7118 2578 -7114
rect 2350 -7166 2578 -7118
rect 2630 -7118 2636 -7114
rect 2852 -7118 2858 -7114
rect 2630 -7166 2858 -7118
rect 2910 -7166 2920 -7114
rect 138 -7800 814 -7748
rect 866 -7800 1094 -7748
rect 1146 -7800 1934 -7748
rect 1986 -7800 2214 -7748
rect 2266 -7800 2276 -7748
rect 2978 -7842 3026 -7010
rect 888 -7894 898 -7842
rect 950 -7894 1178 -7842
rect 1230 -7894 2018 -7842
rect 2070 -7894 2298 -7842
rect 2350 -7894 3026 -7842
rect -390 -8188 210 -8178
rect -390 -8498 210 -8488
rect 3028 -8188 3628 -8178
rect 3028 -8498 3628 -8488
<< via2 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -390 -8488 210 -8188
rect 3028 -8488 3628 -8188
<< metal3 >>
rect -400 1016 220 1021
rect -400 716 -390 1016
rect 210 716 220 1016
rect -400 711 220 716
rect 3018 1016 3638 1021
rect 3018 716 3028 1016
rect 3628 716 3638 1016
rect 3018 711 3638 716
rect -400 -8188 220 -8183
rect -400 -8488 -390 -8188
rect 210 -8488 220 -8188
rect -400 -8493 220 -8488
rect 3018 -8188 3638 -8183
rect 3018 -8488 3028 -8188
rect 3628 -8488 3638 -8188
rect 3018 -8493 3638 -8488
<< via3 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -390 -8488 210 -8188
rect 3028 -8488 3628 -8188
<< metal4 >>
rect -391 1016 211 1017
rect -391 716 -390 1016
rect 210 716 211 1016
rect -391 715 211 716
rect 3027 1016 3629 1017
rect 3027 716 3028 1016
rect 3628 716 3629 1016
rect 3027 715 3629 716
rect -391 -8188 211 -8187
rect -391 -8488 -390 -8188
rect 210 -8488 211 -8188
rect -391 -8489 211 -8488
rect 3027 -8188 3629 -8187
rect 3027 -8488 3028 -8188
rect 3628 -8488 3629 -8188
rect 3027 -8489 3629 -8488
<< labels >>
rlabel metal1 706 670 806 770 1 VDD
port 1 n
rlabel metal1 154 -6156 254 -6056 1 Vioplus
port 6 n
rlabel metal1 2750 -6256 2850 -6156 1 Viominus
port 7 n
rlabel metal1 3274 -1892 3374 -1792 1 CLK
port 3 n
rlabel metal1 3184 -7120 3284 -7020 1 VSS
port 8 n
rlabel metal1 2368 -1448 2468 -1348 1 Voutminus
port 5 n
rlabel metal1 34 -1400 134 -1300 1 Voutplus
port 4 n
<< end >>
