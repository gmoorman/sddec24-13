** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/2stageOpamp.sch
.subckt 2stageOpamp Vinm Vinp Vout VSS VDD Vb1 Vb2 Vb3
*.PININFO Vinm:I Vinp:I Vout:O VSS:I VDD:I Vb1:I Vb2:I Vb3:I
XM8 Vout net1 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=6 nf=1 m=8
XM2 Vout Vb1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=9 nf=1 m=3
XC2 net2 Vout sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=4
XM5 net5 Vb3 net6 VSS sky130_fd_pr__nfet_01v8 L=1 W=4 nf=1 m=3
XM17 net1 Vb3 net7 VSS sky130_fd_pr__nfet_01v8 L=1 W=4 nf=1 m=3
XM3 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=8 nf=1 m=1
XM19 net7 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=8 nf=1 m=1
XM11 net8 Vb1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=9 nf=1 m=2
XM1 net6 Vinm net8 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=3
XM15 net7 Vinp net8 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=3
XM7 net3 Vb1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=9 nf=1 m=1
XM21 net4 Vb1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=9 nf=1 m=1
XM9 net5 Vb2 net3 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=9 nf=1 m=1
XM23 net1 Vb2 net4 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=9 nf=1 m=1
XR1 net2 net1 VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.1 mult=1 m=1
.ends
.end
