* NGSPICE file created from combination_test_WORKING.ext - technology: sky130B

.subckt combination_test_WORKING VDD CLK Voutplus Voutminus Vioplus Viominus VSS
X0 Voutplus.t2 CLK.t0 a_206_n3829.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X1 Voutminus.t0 CLK.t1 a_206_n3009.t0 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X2 a_294_n6912.t0 Viominus.t0 VSS.t6 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X3 Voutminus.t1 CLK.t2 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X4 a_294_n7610# Vioplus.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X5 Voutminus CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15 M=9
X6 a_294_n7610# Vioplus VSS VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15 M=9
X7 Voutminus.t2 Voutplus.t3 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X8 Voutplus.t1 CLK.t3 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X9 a_206_n3829.t0 Voutminus.t3 a_294_n7610# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X10 Voutplus.t0 Voutminus.t4 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X11 Voutplus CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15 M=9
X12 a_206_n3009.t1 Voutplus.t4 a_294_n6912.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X13 Voutminus Voutplus VDD VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X14 Voutplus Voutminus VDD VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
R0 CLK.n19 CLK.n17 566.539
R1 CLK.n10 CLK.n8 566.519
R2 CLK.n2 CLK.n0 566.519
R3 CLK.n35 CLK.n34 565.846
R4 CLK.n33 CLK.n32 565.846
R5 CLK.n31 CLK.n30 565.846
R6 CLK.n29 CLK.n28 565.846
R7 CLK.n27 CLK.n26 565.846
R8 CLK.n25 CLK.n24 565.846
R9 CLK.n23 CLK.n22 565.846
R10 CLK.n21 CLK.n20 565.846
R11 CLK.n19 CLK.n18 565.846
R12 CLK.n10 CLK.n9 565.846
R13 CLK.n12 CLK.n11 565.846
R14 CLK.n14 CLK.n13 565.846
R15 CLK.n15 CLK.t3 565.846
R16 CLK.n7 CLK.t2 565.846
R17 CLK.n6 CLK.n5 565.846
R18 CLK.n4 CLK.n3 565.846
R19 CLK.n2 CLK.n1 565.846
R20 CLK.n56 CLK.n55 551.386
R21 CLK.n54 CLK.n53 551.386
R22 CLK.n52 CLK.n51 551.386
R23 CLK.n50 CLK.n49 551.386
R24 CLK.n48 CLK.n47 551.386
R25 CLK.n46 CLK.n45 551.386
R26 CLK.n44 CLK.n43 551.386
R27 CLK.n42 CLK.t1 551.386
R28 CLK.n41 CLK.n40 551.386
R29 CLK.n39 CLK.n38 551.386
R30 CLK.n58 CLK.n57 551.38
R31 CLK.n60 CLK.n59 551.38
R32 CLK.n62 CLK.n61 551.38
R33 CLK.n64 CLK.n63 551.38
R34 CLK.n66 CLK.n65 551.38
R35 CLK.n68 CLK.n67 551.38
R36 CLK.n69 CLK.t0 551.38
R37 CLK.n71 CLK.n70 551.38
R38 CLK.n73 CLK.n72 551.38
R39 CLK.n75 CLK.n37 542.38
R40 CLK.n76 CLK.n75 10.9256
R41 CLK.n77 CLK.n76 10.0607
R42 CLK.n75 CLK.n74 9.0005
R43 CLK.n36 CLK.n35 6.20021
R44 CLK.n58 CLK.n56 4.52935
R45 CLK.n74 CLK.n39 4.52935
R46 CLK.n36 CLK.n16 3.65435
R47 CLK.n76 CLK.n36 1.23264
R48 CLK.n16 CLK.n7 1.01012
R49 CLK.n16 CLK.n15 1.01012
R50 CLK.n21 CLK.n19 0.693577
R51 CLK.n23 CLK.n21 0.693577
R52 CLK.n25 CLK.n23 0.693577
R53 CLK.n27 CLK.n25 0.693577
R54 CLK.n29 CLK.n27 0.693577
R55 CLK.n31 CLK.n29 0.693577
R56 CLK.n33 CLK.n31 0.693577
R57 CLK.n35 CLK.n33 0.693577
R58 CLK.n41 CLK.n39 0.673577
R59 CLK.n42 CLK.n41 0.673577
R60 CLK.n44 CLK.n42 0.673577
R61 CLK.n46 CLK.n44 0.673577
R62 CLK.n48 CLK.n46 0.673577
R63 CLK.n50 CLK.n48 0.673577
R64 CLK.n52 CLK.n50 0.673577
R65 CLK.n54 CLK.n52 0.673577
R66 CLK.n56 CLK.n54 0.673577
R67 CLK.n74 CLK.n73 0.673577
R68 CLK.n73 CLK.n71 0.673577
R69 CLK.n71 CLK.n69 0.673577
R70 CLK.n69 CLK.n68 0.673577
R71 CLK.n68 CLK.n66 0.673577
R72 CLK.n66 CLK.n64 0.673577
R73 CLK.n64 CLK.n62 0.673577
R74 CLK.n62 CLK.n60 0.673577
R75 CLK.n60 CLK.n58 0.673577
R76 CLK.n4 CLK.n2 0.673577
R77 CLK.n6 CLK.n4 0.673577
R78 CLK.n7 CLK.n6 0.673577
R79 CLK.n15 CLK.n14 0.673577
R80 CLK.n14 CLK.n12 0.673577
R81 CLK.n12 CLK.n10 0.673577
R82 CLK.n77 CLK 0.07175
R83 CLK CLK.n77 0.05425
R84 a_206_n3829.t1 a_206_n3829.t0 107.681
R85 Voutplus.t4 Voutplus.n3 1086.18
R86 Voutplus.n2 Voutplus.n1 582.394
R87 Voutplus.n2 Voutplus.t3 557.25
R88 Voutplus.n4 Voutplus.t4 555.361
R89 Voutplus.n0 Voutplus.t0 124.022
R90 Voutplus.n0 Voutplus.t1 123.349
R91 Voutplus.n4 Voutplus.t2 52.3995
R92 Voutplus.n5 Voutplus.n4 35.4524
R93 Voutplus Voutplus.n0 13.55
R94 Voutplus.n5 Voutplus.n2 5.15969
R95 Voutplus Voutplus.n5 1.44815
R96 VSS.n7 VSS.n6 8103.64
R97 VSS.n9 VSS.n6 8103.64
R98 VSS.n7 VSS.n3 8103.64
R99 VSS.n9 VSS.n3 8103.64
R100 VSS.t3 VSS.n7 928.809
R101 VSS.n9 VSS.t0 826.663
R102 VSS.n10 VSS.n5 674.944
R103 VSS.n11 VSS.n10 674.944
R104 VSS.n11 VSS.n2 674.944
R105 VSS.n5 VSS.n2 674.944
R106 VSS.t0 VSS.t2 357.517
R107 VSS.t4 VSS.t3 178.758
R108 VSS.t5 VSS.t4 178.758
R109 VSS.t2 VSS.n8 140.453
R110 VSS.n14 VSS.t1 53.6536
R111 VSS.n14 VSS.t6 51.4503
R112 VSS.n8 VSS.t5 38.3058
R113 VSS VSS.n14 16.2958
R114 VSS.n11 VSS.n3 10.2637
R115 VSS.n8 VSS.n3 10.2637
R116 VSS.n6 VSS.n5 10.2637
R117 VSS.n8 VSS.n6 10.2637
R118 VSS.n10 VSS.n9 6.29082
R119 VSS.n7 VSS.n2 6.29082
R120 VSS.n4 VSS.n0 5.87885
R121 VSS.n4 VSS.n1 5.87885
R122 VSS.n12 VSS.n1 5.00279
R123 VSS.n13 VSS.n12 3.02064
R124 VSS.n13 VSS.n0 1.98264
R125 VSS VSS.n13 1.59871
R126 VSS.n5 VSS.n4 0.166571
R127 VSS.n12 VSS.n11 0.166571
R128 VSS.n10 VSS.n1 0.11675
R129 VSS.n2 VSS.n0 0.11675
R130 a_206_n3009.t0 a_206_n3009.t1 87.8097
R131 Voutminus.t3 Voutminus.n1 1103.9
R132 Voutminus.n4 Voutminus.n3 572.678
R133 Voutminus.n4 Voutminus.t4 567.236
R134 Voutminus.n2 Voutminus.t3 556.408
R135 Voutminus.n0 Voutminus.t2 124.022
R136 Voutminus.n0 Voutminus.t1 123.349
R137 Voutminus.n2 Voutminus.t0 51.7514
R138 Voutminus.n6 Voutminus.n0 15.3144
R139 Voutminus.n5 Voutminus.n2 10.6996
R140 Voutminus.n6 Voutminus.n5 10.4308
R141 Voutminus.n5 Voutminus.n4 2.9404
R142 Voutminus Voutminus.n6 0.149538
R143 Viominus.n3 Viominus.n1 552.063
R144 Viominus.n7 Viominus.n6 551.39
R145 Viominus.n5 Viominus.n4 551.39
R146 Viominus.n9 Viominus.n8 551.384
R147 Viominus.n11 Viominus.n10 551.384
R148 Viominus.n12 Viominus.t0 551.384
R149 Viominus.n14 Viominus.n13 551.384
R150 Viominus.n16 Viominus.n15 551.384
R151 Viominus.n3 Viominus.n2 551.342
R152 Viominus.n17 Viominus.n0 542.384
R153 Viominus.n17 Viominus.n16 9.67358
R154 Viominus.n9 Viominus.n7 4.81947
R155 Viominus.n5 Viominus.n3 2.01973
R156 Viominus.n16 Viominus.n14 2.01973
R157 Viominus.n12 Viominus.n11 2.01973
R158 Viominus.n7 Viominus.n5 0.673577
R159 Viominus.n14 Viominus.n12 0.673577
R160 Viominus.n11 Viominus.n9 0.673577
R161 Viominus Viominus.n17 0.300274
R162 a_294_n6912.t0 a_294_n6912.t1 131.213
R163 VDD.n7 VDD.n3 3093.63
R164 VDD.n9 VDD.n3 3093.63
R165 VDD.n9 VDD.n6 3093.63
R166 VDD.n7 VDD.n6 3093.63
R167 VDD.t4 VDD.n6 554.597
R168 VDD.t2 VDD.n3 504.228
R169 VDD.n5 VDD.n2 432.257
R170 VDD.n11 VDD.n2 432.257
R171 VDD.n10 VDD.n5 432.257
R172 VDD.n11 VDD.n10 432.257
R173 VDD.n14 VDD.t5 125.6
R174 VDD.n16 VDD.t3 124.927
R175 VDD.n15 VDD.t1 124.927
R176 VDD.n14 VDD.t7 124.927
R177 VDD.t6 VDD.t4 89.2622
R178 VDD.t0 VDD.t2 89.2622
R179 VDD.n8 VDD.t0 69.8159
R180 VDD.n8 VDD.t6 19.4468
R181 VDD VDD.n16 10.164
R182 VDD.n6 VDD.n5 5.0005
R183 VDD.n11 VDD.n3 5.0005
R184 VDD.n12 VDD.n1 3.76278
R185 VDD.n4 VDD.n1 3.76278
R186 VDD.n7 VDD.n2 3.24611
R187 VDD.n8 VDD.n7 3.24611
R188 VDD.n10 VDD.n9 3.24611
R189 VDD.n9 VDD.n8 3.24611
R190 VDD.n4 VDD.n0 2.88671
R191 VDD.n13 VDD.n12 1.92355
R192 VDD.n13 VDD.n0 0.96367
R193 VDD.n15 VDD.n14 0.673577
R194 VDD.n16 VDD.n15 0.673577
R195 VDD VDD.n13 0.591846
R196 VDD.n12 VDD.n11 0.282318
R197 VDD.n5 VDD.n4 0.282318
R198 VDD.n10 VDD.n1 0.166571
R199 VDD.n2 VDD.n0 0.166571
R200 Vioplus.n14 Vioplus.n13 542.548
R201 Vioplus.n11 Vioplus.n10 542.548
R202 Vioplus.n1 Vioplus.t0 542.548
R203 Vioplus.n4 Vioplus.n3 542.548
R204 Vioplus.n14 Vioplus.n12 542.542
R205 Vioplus.n11 Vioplus.n9 542.542
R206 Vioplus.n1 Vioplus.n0 542.542
R207 Vioplus.n4 Vioplus.n2 542.542
R208 Vioplus.n8 Vioplus.n7 542.463
R209 Vioplus.n8 Vioplus.n6 542.458
R210 Vioplus.n17 Vioplus.n16 9.19693
R211 Vioplus.n15 Vioplus.n14 6.48264
R212 Vioplus.n5 Vioplus.n4 5.83979
R213 Vioplus.n16 Vioplus.n15 5.0005
R214 Vioplus.n17 Vioplus.n5 3.46479
R215 Vioplus.n15 Vioplus.n11 1.48264
R216 Vioplus.n16 Vioplus.n8 1.46479
R217 Vioplus.n5 Vioplus.n1 0.839786
R218 Vioplus Vioplus.n17 0.304071
C0 Vioplus Viominus 0.746227f
C1 Vioplus Voutplus 0.007055f
C2 Viominus Voutplus 0.003519f
C3 Vioplus Voutminus 1.64e-19
C4 Viominus Voutminus 0.00352f
C5 CLK Voutplus 5.05098f
C6 Voutplus Voutminus 1.36036f
C7 Voutplus VDD 10.2038f
C8 Vioplus a_294_n7610# 0.74135f
C9 Viominus a_294_n7610# 0.295933f
C10 Voutplus a_294_n7610# 0.066969f
C11 CLK Voutminus 6.14009f
C12 CLK VDD 9.47672f
C13 Voutminus VDD 9.96877f
C14 CLK a_294_n7610# 4.27e-20
C15 Voutminus a_294_n7610# 0.163493f
C16 Vioplus VSS 4.89194f
C17 Viominus VSS 3.243847f
C18 Voutplus VSS 4.459104f
C19 CLK VSS 7.391452f
C20 Voutminus VSS 4.023736f
C21 VDD VSS 48.75097f
C22 a_294_n7610# VSS 8.907901f
C23 VDD.n0 VSS 0.596545f
C24 VDD.n1 VSS 0.575815f
C25 VDD.n2 VSS 0.514341f
C26 VDD.n3 VSS 4.68973f
C27 VDD.n4 VSS 0.924509f
C28 VDD.n5 VSS 0.517698f
C29 VDD.n6 VSS 5.0447f
C30 VDD.t4 VSS 4.53615f
C31 VDD.t6 VSS 0.765055f
C32 VDD.t2 VSS 4.18215f
C33 VDD.t0 VSS 1.11954f
C34 VDD.n7 VSS 0.637232f
C35 VDD.n8 VSS 0.628197f
C36 VDD.n9 VSS 0.637232f
C37 VDD.n10 VSS 0.514341f
C38 VDD.n11 VSS 0.517698f
C39 VDD.n12 VSS 0.69862f
C40 VDD.n13 VSS 0.686525f
C41 VDD.t5 VSS 0.04827f
C42 VDD.t7 VSS 0.044577f
C43 VDD.n14 VSS 0.845197f
C44 VDD.t1 VSS 0.044577f
C45 VDD.n15 VSS 0.159699f
C46 VDD.t3 VSS 0.044577f
C47 VDD.n16 VSS 0.554767f
C48 a_294_n6912.t1 VSS 0.982807f
C49 a_294_n6912.t0 VSS 1.11719f
C50 Viominus.n0 VSS 0.038153f
C51 Viominus.n1 VSS 0.039135f
C52 Viominus.n2 VSS 0.039042f
C53 Viominus.n3 VSS 0.238341f
C54 Viominus.n4 VSS 0.039032f
C55 Viominus.n5 VSS 0.153185f
C56 Viominus.n6 VSS 0.039032f
C57 Viominus.n7 VSS 0.281327f
C58 Viominus.n8 VSS 0.039027f
C59 Viominus.n9 VSS 0.299575f
C60 Viominus.n10 VSS 0.039027f
C61 Viominus.n11 VSS 0.152941f
C62 Viominus.t0 VSS 0.039027f
C63 Viominus.n12 VSS 0.152941f
C64 Viominus.n13 VSS 0.039027f
C65 Viominus.n14 VSS 0.152941f
C66 Viominus.n15 VSS 0.039027f
C67 Viominus.n16 VSS 0.182268f
C68 Viominus.n17 VSS 0.057204f
C69 Voutminus.t2 VSS 0.373067f
C70 Voutminus.t1 VSS 0.36727f
C71 Voutminus.n0 VSS 4.95382f
C72 Voutminus.n1 VSS 0.521294f
C73 Voutminus.t3 VSS 0.551459f
C74 Voutminus.t0 VSS 0.404434f
C75 Voutminus.n2 VSS 5.22831f
C76 Voutminus.t4 VSS 0.297302f
C77 Voutminus.n3 VSS 0.310636f
C78 Voutminus.n4 VSS 3.30533f
C79 Voutminus.n5 VSS 4.95304f
C80 Voutminus.n6 VSS 1.70453f
C81 a_206_n3009.t1 VSS 5.25228f
C82 a_206_n3009.t0 VSS 5.34772f
C83 Voutplus.t0 VSS 0.421038f
C84 Voutplus.t1 VSS 0.414495f
C85 Voutplus.n0 VSS 5.38868f
C86 Voutplus.t3 VSS 0.329803f
C87 Voutplus.n1 VSS 0.396193f
C88 Voutplus.n2 VSS 3.42741f
C89 Voutplus.t2 VSS 0.485682f
C90 Voutplus.n3 VSS 0.47775f
C91 Voutplus.t4 VSS 0.508627f
C92 Voutplus.n4 VSS 6.54139f
C93 Voutplus.n5 VSS 1.48899f
C94 a_206_n3829.t0 VSS 3.26775f
C95 a_206_n3829.t1 VSS 3.03225f
C96 CLK.n0 VSS 0.207276f
C97 CLK.n1 VSS 0.206996f
C98 CLK.n2 VSS 0.522139f
C99 CLK.n3 VSS 0.206996f
C100 CLK.n4 VSS 0.287044f
C101 CLK.n5 VSS 0.206996f
C102 CLK.n6 VSS 0.287044f
C103 CLK.t2 VSS 0.206996f
C104 CLK.n7 VSS 0.321822f
C105 CLK.n8 VSS 0.207276f
C106 CLK.n9 VSS 0.206996f
C107 CLK.n10 VSS 0.522139f
C108 CLK.n11 VSS 0.206996f
C109 CLK.n12 VSS 0.287044f
C110 CLK.n13 VSS 0.206996f
C111 CLK.n14 VSS 0.287044f
C112 CLK.t3 VSS 0.206996f
C113 CLK.n15 VSS 0.321822f
C114 CLK.n16 VSS 0.597953f
C115 CLK.n17 VSS 0.207282f
C116 CLK.n18 VSS 0.206996f
C117 CLK.n19 VSS 0.516171f
C118 CLK.n20 VSS 0.206996f
C119 CLK.n21 VSS 0.28307f
C120 CLK.n22 VSS 0.206996f
C121 CLK.n23 VSS 0.28307f
C122 CLK.n24 VSS 0.206996f
C123 CLK.n25 VSS 0.28307f
C124 CLK.n26 VSS 0.206996f
C125 CLK.n27 VSS 0.28307f
C126 CLK.n28 VSS 0.206996f
C127 CLK.n29 VSS 0.28307f
C128 CLK.n30 VSS 0.206996f
C129 CLK.n31 VSS 0.28307f
C130 CLK.n32 VSS 0.206996f
C131 CLK.n33 VSS 0.28307f
C132 CLK.n34 VSS 0.206996f
C133 CLK.n35 VSS 0.851343f
C134 CLK.n36 VSS 1.19268f
C135 CLK.n37 VSS 0.200931f
C136 CLK.n38 VSS 0.20405f
C137 CLK.n39 VSS 0.696894f
C138 CLK.n40 VSS 0.20405f
C139 CLK.n41 VSS 0.285519f
C140 CLK.t1 VSS 0.20405f
C141 CLK.n42 VSS 0.285519f
C142 CLK.n43 VSS 0.20405f
C143 CLK.n44 VSS 0.285519f
C144 CLK.n45 VSS 0.20405f
C145 CLK.n46 VSS 0.285519f
C146 CLK.n47 VSS 0.20405f
C147 CLK.n48 VSS 0.285519f
C148 CLK.n49 VSS 0.20405f
C149 CLK.n50 VSS 0.285519f
C150 CLK.n51 VSS 0.20405f
C151 CLK.n52 VSS 0.285519f
C152 CLK.n53 VSS 0.20405f
C153 CLK.n54 VSS 0.285519f
C154 CLK.n55 VSS 0.20405f
C155 CLK.n56 VSS 0.696894f
C156 CLK.n57 VSS 0.203349f
C157 CLK.n58 VSS 0.696219f
C158 CLK.n59 VSS 0.203349f
C159 CLK.n60 VSS 0.284844f
C160 CLK.n61 VSS 0.203349f
C161 CLK.n62 VSS 0.284844f
C162 CLK.n63 VSS 0.203349f
C163 CLK.n64 VSS 0.284844f
C164 CLK.n65 VSS 0.203349f
C165 CLK.n66 VSS 0.284844f
C166 CLK.n67 VSS 0.203349f
C167 CLK.n68 VSS 0.284844f
C168 CLK.t0 VSS 0.203349f
C169 CLK.n69 VSS 0.284844f
C170 CLK.n70 VSS 0.203349f
C171 CLK.n71 VSS 0.284844f
C172 CLK.n72 VSS 0.203349f
C173 CLK.n73 VSS 0.284844f
C174 CLK.n74 VSS 0.550488f
C175 CLK.n75 VSS 0.264976f
C176 CLK.n76 VSS 0.413662f
C177 CLK.n77 VSS 0.182118f
.ends

