** sch_path: /home/jaxie963/caravel_pls_man_analog/caravel_user_project_analog/xschem/Preamp_noBias.sch
.subckt Preamp_noBias VDD VSS Vinplus Vinminus Vioplus Viominus i_in
*.PININFO VDD:B VSS:B Vinplus:B Vinminus:B Vioplus:B Viominus:B i_in:B
XM11 Viominus Vinminus net1 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=4
XM12 Vioplus Vinplus net1 VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=4
XM14 net1 i_in VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=10
XR2 VSS Vioplus VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.751 mult=1 m=1
XR1 Viominus VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.751 mult=1 m=1
.ends
.end
