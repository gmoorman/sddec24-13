magic
tech sky130B
timestamp 1730400109
<< checkpaint >>
rect -630 -330 1870 2135
rect -630 -1830 730 -330
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
use 1T1Rcomp  x1 ~/reram/caravel_user_project_analog/mag
timestamp 1730396854
transform 1 0 90 0 1 90
box -90 210 220 1415
use 1T1Rcomp  x2
timestamp 1730396854
transform 1 0 400 0 1 90
box -90 210 220 1415
use 1T1Rcomp  x3
timestamp 1730396854
transform 1 0 710 0 1 90
box -90 210 220 1415
use 1T1Rcomp  x4
timestamp 1730396854
transform 1 0 1020 0 1 90
box -90 210 220 1415
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 BL2
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 BL1
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 VSS
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 WL1
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 WL2
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 SL1
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 SL2
port 6 nsew
<< end >>
