magic
tech sky130B
magscale 1 2
timestamp 1733718626
<< viali >>
rect 3985 5321 4019 5355
rect 4353 5321 4387 5355
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 3157 5185 3191 5219
rect 3433 5185 3467 5219
rect 3801 5185 3835 5219
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 4537 5185 4571 5219
rect 4813 5185 4847 5219
rect 4997 5185 5031 5219
rect 5273 5185 5307 5219
rect 5549 5185 5583 5219
rect 5733 5185 5767 5219
rect 5917 5185 5951 5219
rect 6009 5185 6043 5219
rect 1593 5117 1627 5151
rect 4169 5117 4203 5151
rect 5457 5117 5491 5151
rect 3341 5049 3375 5083
rect 5365 5049 5399 5083
rect 3065 4981 3099 5015
rect 3617 4981 3651 5015
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 6193 4981 6227 5015
rect 3065 4777 3099 4811
rect 5365 4777 5399 4811
rect 5733 4777 5767 4811
rect 3617 4709 3651 4743
rect 2145 4641 2179 4675
rect 2605 4573 2639 4607
rect 2881 4573 2915 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 4905 4573 4939 4607
rect 4997 4573 5031 4607
rect 5365 4573 5399 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6009 4573 6043 4607
rect 6101 4573 6135 4607
rect 6193 4573 6227 4607
rect 4077 4505 4111 4539
rect 3341 4437 3375 4471
rect 4813 4437 4847 4471
rect 5181 4437 5215 4471
rect 4721 4233 4755 4267
rect 4537 4165 4571 4199
rect 5457 4165 5491 4199
rect 3709 4097 3743 4131
rect 4261 4097 4295 4131
rect 4353 4097 4387 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 4905 4097 4939 4131
rect 5174 4097 5208 4131
rect 5365 4097 5399 4131
rect 5641 4097 5675 4131
rect 5917 4097 5951 4131
rect 6101 4097 6135 4131
rect 3893 3893 3927 3927
rect 3985 3893 4019 3927
rect 4169 3893 4203 3927
rect 4261 3689 4295 3723
rect 5181 3689 5215 3723
rect 5917 3689 5951 3723
rect 6009 3689 6043 3723
rect 6469 3689 6503 3723
rect 2789 3485 2823 3519
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 4813 3485 4847 3519
rect 4905 3485 4939 3519
rect 4997 3485 5031 3519
rect 5273 3485 5307 3519
rect 5457 3485 5491 3519
rect 5733 3485 5767 3519
rect 6193 3485 6227 3519
rect 6285 3485 6319 3519
rect 1593 3417 1627 3451
rect 6009 3417 6043 3451
rect 3985 3349 4019 3383
rect 4353 3349 4387 3383
rect 5457 3145 5491 3179
rect 4629 3077 4663 3111
rect 5181 3077 5215 3111
rect 5365 3077 5399 3111
rect 4261 3009 4295 3043
rect 4537 3009 4571 3043
rect 4813 3009 4847 3043
rect 5089 3009 5123 3043
rect 5641 3009 5675 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 5292 2941 5326 2975
rect 4997 2873 5031 2907
rect 4445 2805 4479 2839
rect 4905 2601 4939 2635
rect 5641 2601 5675 2635
rect 5365 2465 5399 2499
rect 2697 2397 2731 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 5273 2397 5307 2431
rect 5457 2397 5491 2431
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 1593 2329 1627 2363
rect 4997 2261 5031 2295
rect 6009 2261 6043 2295
<< metal1 >>
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3016 5868 6592 5896
rect 3016 5856 3022 5868
rect 6564 5840 6592 5868
rect 6546 5788 6552 5840
rect 6604 5788 6610 5840
rect 3326 5720 3332 5772
rect 3384 5760 3390 5772
rect 3384 5732 7052 5760
rect 3384 5720 3390 5732
rect 7024 5704 7052 5732
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5626 5692 5632 5704
rect 4212 5664 5632 5692
rect 4212 5652 4218 5664
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 3660 5596 6408 5624
rect 3660 5584 3666 5596
rect 6380 5568 6408 5596
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 5718 5556 5724 5568
rect 3752 5528 5724 5556
rect 3752 5516 3758 5528
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6362 5516 6368 5568
rect 6420 5516 6426 5568
rect 1104 5466 6968 5488
rect 1104 5414 2376 5466
rect 2428 5414 2440 5466
rect 2492 5414 2504 5466
rect 2556 5414 2568 5466
rect 2620 5414 2632 5466
rect 2684 5414 3802 5466
rect 3854 5414 3866 5466
rect 3918 5414 3930 5466
rect 3982 5414 3994 5466
rect 4046 5414 4058 5466
rect 4110 5414 5228 5466
rect 5280 5414 5292 5466
rect 5344 5414 5356 5466
rect 5408 5414 5420 5466
rect 5472 5414 5484 5466
rect 5536 5414 6654 5466
rect 6706 5414 6718 5466
rect 6770 5414 6782 5466
rect 6834 5414 6846 5466
rect 6898 5414 6910 5466
rect 6962 5414 6968 5466
rect 1104 5392 6968 5414
rect 3510 5352 3516 5364
rect 2884 5324 3516 5352
rect 2682 5176 2688 5228
rect 2740 5176 2746 5228
rect 2884 5225 2912 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3844 5324 3985 5352
rect 3844 5312 3850 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 4338 5312 4344 5364
rect 4396 5312 4402 5364
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 5902 5352 5908 5364
rect 4488 5324 5908 5352
rect 4488 5312 4494 5324
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 2976 5256 4200 5284
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 992 5120 1593 5148
rect 992 5108 998 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 2976 5080 3004 5256
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3160 5148 3188 5179
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3384 5188 3433 5216
rect 3384 5176 3390 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3660 5188 3801 5216
rect 3660 5176 3666 5188
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 4028 5188 4077 5216
rect 4028 5176 4034 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 3528 5148 3556 5176
rect 4172 5157 4200 5256
rect 4448 5256 5120 5284
rect 4249 5220 4307 5225
rect 4249 5219 4378 5220
rect 4249 5185 4261 5219
rect 4295 5216 4378 5219
rect 4448 5216 4476 5256
rect 4295 5192 4476 5216
rect 4295 5185 4307 5192
rect 4350 5188 4476 5192
rect 4249 5179 4307 5185
rect 3160 5120 3556 5148
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5117 4215 5151
rect 4448 5148 4476 5188
rect 4522 5176 4528 5228
rect 4580 5176 4586 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4816 5148 4844 5179
rect 4982 5176 4988 5228
rect 5040 5176 5046 5228
rect 5092 5216 5120 5256
rect 5166 5244 5172 5296
rect 5224 5284 5230 5296
rect 5224 5256 6040 5284
rect 5224 5244 5230 5256
rect 5092 5188 5212 5216
rect 5074 5148 5080 5160
rect 4448 5120 4660 5148
rect 4816 5120 5080 5148
rect 4157 5111 4215 5117
rect 2924 5052 3004 5080
rect 3329 5083 3387 5089
rect 2924 5040 2930 5052
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 4338 5080 4344 5092
rect 3375 5052 4344 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 4338 5040 4344 5052
rect 4396 5080 4402 5092
rect 4522 5080 4528 5092
rect 4396 5052 4528 5080
rect 4396 5040 4402 5052
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 3510 5012 3516 5024
rect 3099 4984 3516 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4154 5012 4160 5024
rect 3651 4984 4160 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4632 5012 4660 5120
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5184 5148 5212 5188
rect 5258 5176 5264 5228
rect 5316 5176 5322 5228
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 5902 5176 5908 5228
rect 5960 5176 5966 5228
rect 6012 5225 6040 5256
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 5368 5148 5396 5176
rect 5184 5120 5396 5148
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5491 5120 5948 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 4890 5040 4896 5092
rect 4948 5080 4954 5092
rect 5353 5083 5411 5089
rect 5353 5080 5365 5083
rect 4948 5052 5365 5080
rect 4948 5040 4954 5052
rect 5353 5049 5365 5052
rect 5399 5049 5411 5083
rect 5920 5080 5948 5120
rect 6454 5080 6460 5092
rect 5920 5052 6460 5080
rect 5353 5043 5411 5049
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 4304 4984 4660 5012
rect 4304 4972 4310 4984
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 5040 4984 5089 5012
rect 5040 4972 5046 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5077 4975 5135 4981
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5500 4984 5733 5012
rect 5500 4972 5506 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6270 5012 6276 5024
rect 6227 4984 6276 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 1104 4922 6808 4944
rect 1104 4870 1663 4922
rect 1715 4870 1727 4922
rect 1779 4870 1791 4922
rect 1843 4870 1855 4922
rect 1907 4870 1919 4922
rect 1971 4870 3089 4922
rect 3141 4870 3153 4922
rect 3205 4870 3217 4922
rect 3269 4870 3281 4922
rect 3333 4870 3345 4922
rect 3397 4870 4515 4922
rect 4567 4870 4579 4922
rect 4631 4870 4643 4922
rect 4695 4870 4707 4922
rect 4759 4870 4771 4922
rect 4823 4870 5941 4922
rect 5993 4870 6005 4922
rect 6057 4870 6069 4922
rect 6121 4870 6133 4922
rect 6185 4870 6197 4922
rect 6249 4870 6808 4922
rect 1104 4848 6808 4870
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3970 4808 3976 4820
rect 3099 4780 3976 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4062 4768 4068 4820
rect 4120 4768 4126 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4706 4808 4712 4820
rect 4212 4780 4712 4808
rect 4212 4768 4218 4780
rect 4706 4768 4712 4780
rect 4764 4808 4770 4820
rect 5166 4808 5172 4820
rect 4764 4780 5172 4808
rect 4764 4768 4770 4780
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5408 4780 5672 4808
rect 5408 4768 5414 4780
rect 3326 4740 3332 4752
rect 2884 4712 3332 4740
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2774 4672 2780 4684
rect 2179 4644 2780 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 2590 4564 2596 4616
rect 2648 4564 2654 4616
rect 2884 4613 2912 4712
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 3602 4700 3608 4752
rect 3660 4700 3666 4752
rect 4080 4740 4108 4768
rect 5442 4740 5448 4752
rect 4080 4712 4292 4740
rect 2958 4632 2964 4684
rect 3016 4632 3022 4684
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2976 4604 3004 4632
rect 3145 4607 3203 4613
rect 3145 4604 3157 4607
rect 2976 4576 3157 4604
rect 2869 4567 2927 4573
rect 3145 4573 3157 4576
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3418 4564 3424 4616
rect 3476 4564 3482 4616
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4264 4613 4292 4712
rect 4632 4712 5448 4740
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3752 4576 3801 4604
rect 3752 4564 3758 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4430 4564 4436 4616
rect 4488 4564 4494 4616
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 4065 4539 4123 4545
rect 4065 4536 4077 4539
rect 2832 4508 4077 4536
rect 2832 4496 2838 4508
rect 4065 4505 4077 4508
rect 4111 4505 4123 4539
rect 4356 4536 4384 4564
rect 4632 4536 4660 4712
rect 5442 4700 5448 4712
rect 5500 4700 5506 4752
rect 5644 4740 5672 4780
rect 5718 4768 5724 4820
rect 5776 4768 5782 4820
rect 5994 4740 6000 4752
rect 5644 4712 6000 4740
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 5644 4644 6224 4672
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4600 5043 4607
rect 5353 4607 5411 4613
rect 5031 4573 5323 4600
rect 4985 4572 5323 4573
rect 4985 4567 5043 4572
rect 4908 4536 4936 4567
rect 4356 4508 4936 4536
rect 4065 4499 4123 4505
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 4522 4468 4528 4480
rect 3375 4440 4528 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 4801 4471 4859 4477
rect 4801 4468 4813 4471
rect 4672 4440 4813 4468
rect 4672 4428 4678 4440
rect 4801 4437 4813 4440
rect 4847 4437 4859 4471
rect 4801 4431 4859 4437
rect 5166 4428 5172 4480
rect 5224 4428 5230 4480
rect 5295 4468 5323 4572
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5552 4604 5580 4632
rect 5644 4613 5672 4644
rect 5399 4576 5580 4604
rect 5629 4607 5687 4613
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 5736 4536 5764 4564
rect 6012 4536 6040 4567
rect 6086 4564 6092 4616
rect 6144 4564 6150 4616
rect 6196 4613 6224 4644
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6270 4604 6276 4616
rect 6227 4576 6276 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 5736 4508 6040 4536
rect 6104 4468 6132 4564
rect 5295 4440 6132 4468
rect 1104 4378 6968 4400
rect 1104 4326 2376 4378
rect 2428 4326 2440 4378
rect 2492 4326 2504 4378
rect 2556 4326 2568 4378
rect 2620 4326 2632 4378
rect 2684 4326 3802 4378
rect 3854 4326 3866 4378
rect 3918 4326 3930 4378
rect 3982 4326 3994 4378
rect 4046 4326 4058 4378
rect 4110 4326 5228 4378
rect 5280 4326 5292 4378
rect 5344 4326 5356 4378
rect 5408 4326 5420 4378
rect 5472 4326 5484 4378
rect 5536 4326 6654 4378
rect 6706 4326 6718 4378
rect 6770 4326 6782 4378
rect 6834 4326 6846 4378
rect 6898 4326 6910 4378
rect 6962 4326 6968 4378
rect 1104 4304 6968 4326
rect 4430 4224 4436 4276
rect 4488 4224 4494 4276
rect 4709 4267 4767 4273
rect 4709 4233 4721 4267
rect 4755 4264 4767 4267
rect 4890 4264 4896 4276
rect 4755 4236 4896 4264
rect 4755 4233 4767 4236
rect 4709 4227 4767 4233
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 6086 4264 6092 4276
rect 5000 4236 6092 4264
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 4448 4196 4476 4224
rect 3568 4168 4476 4196
rect 4525 4199 4583 4205
rect 3568 4156 3574 4168
rect 4264 4137 4292 4168
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 5000 4196 5028 4236
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 5445 4199 5503 4205
rect 5445 4196 5457 4199
rect 4571 4168 5028 4196
rect 5295 4168 5457 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 5295 4152 5323 4168
rect 5445 4165 5457 4168
rect 5491 4165 5503 4199
rect 5445 4159 5503 4165
rect 5276 4150 5323 4152
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 3712 4060 3740 4091
rect 4338 4088 4344 4140
rect 4396 4088 4402 4140
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4798 4128 4804 4140
rect 4663 4100 4804 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4154 4060 4160 4072
rect 3712 4032 4160 4060
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4448 4060 4476 4091
rect 4798 4088 4804 4100
rect 4856 4128 4862 4140
rect 5184 4137 5323 4150
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4856 4100 4905 4128
rect 4856 4088 4862 4100
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 5162 4131 5323 4137
rect 5162 4097 5174 4131
rect 5208 4124 5323 4131
rect 5353 4131 5411 4137
rect 5208 4122 5304 4124
rect 5208 4097 5220 4122
rect 5162 4091 5220 4097
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 4522 4060 4528 4072
rect 4448 4032 4528 4060
rect 4522 4020 4528 4032
rect 4580 4060 4586 4072
rect 5074 4060 5080 4072
rect 4580 4032 5080 4060
rect 4580 4020 4586 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 5380 4060 5408 4091
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5868 4100 5917 4128
rect 5868 4088 5874 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 6052 4100 6101 4128
rect 6052 4088 6058 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 5132 4032 5408 4060
rect 5132 4020 5138 4032
rect 3712 3964 4200 3992
rect 3712 3936 3740 3964
rect 3694 3884 3700 3936
rect 3752 3884 3758 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4172 3933 4200 3964
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 6454 3992 6460 4004
rect 5684 3964 6460 3992
rect 5684 3952 5690 3964
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3893 4215 3927
rect 4157 3887 4215 3893
rect 1104 3834 6808 3856
rect 1104 3782 1663 3834
rect 1715 3782 1727 3834
rect 1779 3782 1791 3834
rect 1843 3782 1855 3834
rect 1907 3782 1919 3834
rect 1971 3782 3089 3834
rect 3141 3782 3153 3834
rect 3205 3782 3217 3834
rect 3269 3782 3281 3834
rect 3333 3782 3345 3834
rect 3397 3782 4515 3834
rect 4567 3782 4579 3834
rect 4631 3782 4643 3834
rect 4695 3782 4707 3834
rect 4759 3782 4771 3834
rect 4823 3782 5941 3834
rect 5993 3782 6005 3834
rect 6057 3782 6069 3834
rect 6121 3782 6133 3834
rect 6185 3782 6197 3834
rect 6249 3782 6808 3834
rect 1104 3760 6808 3782
rect 3970 3720 3976 3732
rect 2792 3692 3976 3720
rect 2792 3525 2820 3692
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 4706 3720 4712 3732
rect 4295 3692 4712 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5626 3720 5632 3732
rect 5215 3692 5632 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5868 3692 5917 3720
rect 5868 3680 5874 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 5994 3680 6000 3732
rect 6052 3680 6058 3732
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6457 3723 6515 3729
rect 6457 3720 6469 3723
rect 6328 3692 6469 3720
rect 6328 3680 6334 3692
rect 6457 3689 6469 3692
rect 6503 3689 6515 3723
rect 6457 3683 6515 3689
rect 4890 3652 4896 3664
rect 3804 3624 4896 3652
rect 3804 3525 3832 3624
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 5718 3652 5724 3664
rect 5295 3624 5724 3652
rect 3878 3544 3884 3596
rect 3936 3544 3942 3596
rect 4430 3584 4436 3596
rect 4080 3556 4436 3584
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1581 3451 1639 3457
rect 1581 3448 1593 3451
rect 992 3420 1593 3448
rect 992 3408 998 3420
rect 1581 3417 1593 3420
rect 1627 3417 1639 3451
rect 3896 3448 3924 3544
rect 4080 3525 4108 3556
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 5295 3584 5323 3624
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 4724 3556 5323 3584
rect 5368 3556 6316 3584
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4212 3488 4537 3516
rect 4212 3476 4218 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 4724 3525 4752 3556
rect 5368 3528 5396 3556
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4672 3488 4721 3516
rect 4672 3476 4678 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5074 3516 5080 3528
rect 5031 3488 5080 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 4908 3448 4936 3479
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5184 3488 5273 3516
rect 5184 3448 5212 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 3896 3420 5212 3448
rect 1581 3411 1639 3417
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4154 3380 4160 3392
rect 4019 3352 4160 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 4341 3383 4399 3389
rect 4341 3380 4353 3383
rect 4304 3352 4353 3380
rect 4304 3340 4310 3352
rect 4341 3349 4353 3352
rect 4387 3349 4399 3383
rect 5276 3380 5304 3479
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5534 3516 5540 3528
rect 5491 3488 5540 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5736 3525 5764 3556
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6288 3525 6316 3556
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 6144 3488 6193 3516
rect 6144 3476 6150 3488
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3417 6055 3451
rect 5997 3411 6055 3417
rect 6012 3380 6040 3411
rect 5276 3352 6040 3380
rect 4341 3343 4399 3349
rect 1104 3290 6968 3312
rect 1104 3238 2376 3290
rect 2428 3238 2440 3290
rect 2492 3238 2504 3290
rect 2556 3238 2568 3290
rect 2620 3238 2632 3290
rect 2684 3238 3802 3290
rect 3854 3238 3866 3290
rect 3918 3238 3930 3290
rect 3982 3238 3994 3290
rect 4046 3238 4058 3290
rect 4110 3238 5228 3290
rect 5280 3238 5292 3290
rect 5344 3238 5356 3290
rect 5408 3238 5420 3290
rect 5472 3238 5484 3290
rect 5536 3238 6654 3290
rect 6706 3238 6718 3290
rect 6770 3238 6782 3290
rect 6834 3238 6846 3290
rect 6898 3238 6910 3290
rect 6962 3238 6968 3290
rect 1104 3216 6968 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 4522 3176 4528 3188
rect 2924 3148 4528 3176
rect 2924 3136 2930 3148
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5445 3179 5503 3185
rect 4764 3148 5304 3176
rect 4764 3136 4770 3148
rect 5276 3120 5304 3148
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 5626 3176 5632 3188
rect 5491 3148 5632 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 4617 3111 4675 3117
rect 4617 3077 4629 3111
rect 4663 3108 4675 3111
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 4663 3080 5181 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 5169 3077 5181 3080
rect 5215 3077 5227 3111
rect 5169 3071 5227 3077
rect 5258 3068 5264 3120
rect 5316 3068 5322 3120
rect 5350 3068 5356 3120
rect 5408 3068 5414 3120
rect 5994 3108 6000 3120
rect 5644 3080 6000 3108
rect 4246 3000 4252 3052
rect 4304 3000 4310 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 4847 3012 4936 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 4540 2836 4568 3003
rect 4798 2836 4804 2848
rect 4479 2808 4804 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 4908 2836 4936 3012
rect 4982 3000 4988 3052
rect 5040 3000 5046 3052
rect 5074 3000 5080 3052
rect 5132 3000 5138 3052
rect 5276 3040 5304 3068
rect 5644 3049 5672 3080
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5276 3012 5641 3040
rect 5629 3009 5641 3012
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 5000 2972 5028 3000
rect 5280 2975 5338 2981
rect 5000 2944 5120 2972
rect 4985 2907 5043 2913
rect 4985 2873 4997 2907
rect 5031 2904 5043 2907
rect 5092 2904 5120 2944
rect 5280 2941 5292 2975
rect 5326 2972 5338 2975
rect 5920 2972 5948 3003
rect 6086 3000 6092 3052
rect 6144 3000 6150 3052
rect 5326 2944 5948 2972
rect 5326 2941 5338 2944
rect 5280 2935 5338 2941
rect 5031 2876 5120 2904
rect 5031 2873 5043 2876
rect 4985 2867 5043 2873
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6104 2904 6132 3000
rect 6362 2932 6368 2984
rect 6420 2932 6426 2984
rect 5868 2876 6132 2904
rect 5868 2864 5874 2876
rect 6380 2836 6408 2932
rect 4908 2808 6408 2836
rect 1104 2746 6808 2768
rect 1104 2694 1663 2746
rect 1715 2694 1727 2746
rect 1779 2694 1791 2746
rect 1843 2694 1855 2746
rect 1907 2694 1919 2746
rect 1971 2694 3089 2746
rect 3141 2694 3153 2746
rect 3205 2694 3217 2746
rect 3269 2694 3281 2746
rect 3333 2694 3345 2746
rect 3397 2694 4515 2746
rect 4567 2694 4579 2746
rect 4631 2694 4643 2746
rect 4695 2694 4707 2746
rect 4759 2694 4771 2746
rect 4823 2694 5941 2746
rect 5993 2694 6005 2746
rect 6057 2694 6069 2746
rect 6121 2694 6133 2746
rect 6185 2694 6197 2746
rect 6249 2694 6808 2746
rect 1104 2672 6808 2694
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5074 2632 5080 2644
rect 4939 2604 5080 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5626 2592 5632 2644
rect 5684 2592 5690 2644
rect 5092 2536 6224 2564
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2774 2428 2780 2440
rect 2731 2400 2780 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5092 2428 5120 2536
rect 6196 2508 6224 2536
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2496 5411 2499
rect 5399 2468 5856 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 4755 2400 5120 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5166 2388 5172 2440
rect 5224 2388 5230 2440
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5828 2437 5856 2468
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 1578 2320 1584 2372
rect 1636 2320 1642 2372
rect 5350 2360 5356 2372
rect 5000 2332 5356 2360
rect 5000 2301 5028 2332
rect 5350 2320 5356 2332
rect 5408 2360 5414 2372
rect 5552 2360 5580 2391
rect 5408 2332 5580 2360
rect 5408 2320 5414 2332
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2261 5043 2295
rect 4985 2255 5043 2261
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 5132 2264 6009 2292
rect 5132 2252 5138 2264
rect 5997 2261 6009 2264
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 1104 2202 6968 2224
rect 1104 2150 2376 2202
rect 2428 2150 2440 2202
rect 2492 2150 2504 2202
rect 2556 2150 2568 2202
rect 2620 2150 2632 2202
rect 2684 2150 3802 2202
rect 3854 2150 3866 2202
rect 3918 2150 3930 2202
rect 3982 2150 3994 2202
rect 4046 2150 4058 2202
rect 4110 2150 5228 2202
rect 5280 2150 5292 2202
rect 5344 2150 5356 2202
rect 5408 2150 5420 2202
rect 5472 2150 5484 2202
rect 5536 2150 6654 2202
rect 6706 2150 6718 2202
rect 6770 2150 6782 2202
rect 6834 2150 6846 2202
rect 6898 2150 6910 2202
rect 6962 2150 6968 2202
rect 1104 2128 6968 2150
rect 4154 2048 4160 2100
rect 4212 2088 4218 2100
rect 5810 2088 5816 2100
rect 4212 2060 5816 2088
rect 4212 2048 4218 2060
rect 5810 2048 5816 2060
rect 5868 2048 5874 2100
<< via1 >>
rect 2964 5856 3016 5908
rect 6552 5788 6604 5840
rect 3332 5720 3384 5772
rect 4160 5652 4212 5704
rect 5632 5652 5684 5704
rect 7012 5652 7064 5704
rect 3608 5584 3660 5636
rect 3700 5516 3752 5568
rect 5724 5516 5776 5568
rect 6368 5516 6420 5568
rect 2376 5414 2428 5466
rect 2440 5414 2492 5466
rect 2504 5414 2556 5466
rect 2568 5414 2620 5466
rect 2632 5414 2684 5466
rect 3802 5414 3854 5466
rect 3866 5414 3918 5466
rect 3930 5414 3982 5466
rect 3994 5414 4046 5466
rect 4058 5414 4110 5466
rect 5228 5414 5280 5466
rect 5292 5414 5344 5466
rect 5356 5414 5408 5466
rect 5420 5414 5472 5466
rect 5484 5414 5536 5466
rect 6654 5414 6706 5466
rect 6718 5414 6770 5466
rect 6782 5414 6834 5466
rect 6846 5414 6898 5466
rect 6910 5414 6962 5466
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 3516 5312 3568 5364
rect 3792 5312 3844 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 4436 5312 4488 5364
rect 5908 5312 5960 5364
rect 940 5108 992 5160
rect 2872 5040 2924 5092
rect 3332 5176 3384 5228
rect 3516 5176 3568 5228
rect 3608 5176 3660 5228
rect 3976 5176 4028 5228
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 5172 5244 5224 5296
rect 4344 5040 4396 5092
rect 4528 5040 4580 5092
rect 3516 4972 3568 5024
rect 4160 4972 4212 5024
rect 4252 4972 4304 5024
rect 5080 5108 5132 5160
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5356 5176 5408 5228
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 4896 5040 4948 5092
rect 6460 5040 6512 5092
rect 4988 4972 5040 5024
rect 5448 4972 5500 5024
rect 6276 4972 6328 5024
rect 1663 4870 1715 4922
rect 1727 4870 1779 4922
rect 1791 4870 1843 4922
rect 1855 4870 1907 4922
rect 1919 4870 1971 4922
rect 3089 4870 3141 4922
rect 3153 4870 3205 4922
rect 3217 4870 3269 4922
rect 3281 4870 3333 4922
rect 3345 4870 3397 4922
rect 4515 4870 4567 4922
rect 4579 4870 4631 4922
rect 4643 4870 4695 4922
rect 4707 4870 4759 4922
rect 4771 4870 4823 4922
rect 5941 4870 5993 4922
rect 6005 4870 6057 4922
rect 6069 4870 6121 4922
rect 6133 4870 6185 4922
rect 6197 4870 6249 4922
rect 3976 4768 4028 4820
rect 4068 4768 4120 4820
rect 4160 4768 4212 4820
rect 4712 4768 4764 4820
rect 5172 4768 5224 4820
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 2780 4632 2832 4684
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 3332 4700 3384 4752
rect 3608 4743 3660 4752
rect 3608 4709 3617 4743
rect 3617 4709 3651 4743
rect 3651 4709 3660 4743
rect 3608 4700 3660 4709
rect 2964 4632 3016 4684
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 3700 4564 3752 4616
rect 4344 4564 4396 4616
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 2780 4496 2832 4548
rect 5448 4700 5500 4752
rect 5724 4811 5776 4820
rect 5724 4777 5733 4811
rect 5733 4777 5767 4811
rect 5767 4777 5776 4811
rect 5724 4768 5776 4777
rect 6000 4700 6052 4752
rect 5540 4632 5592 4684
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 4528 4428 4580 4480
rect 4620 4428 4672 4480
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 5724 4564 5776 4616
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 6276 4564 6328 4616
rect 2376 4326 2428 4378
rect 2440 4326 2492 4378
rect 2504 4326 2556 4378
rect 2568 4326 2620 4378
rect 2632 4326 2684 4378
rect 3802 4326 3854 4378
rect 3866 4326 3918 4378
rect 3930 4326 3982 4378
rect 3994 4326 4046 4378
rect 4058 4326 4110 4378
rect 5228 4326 5280 4378
rect 5292 4326 5344 4378
rect 5356 4326 5408 4378
rect 5420 4326 5472 4378
rect 5484 4326 5536 4378
rect 6654 4326 6706 4378
rect 6718 4326 6770 4378
rect 6782 4326 6834 4378
rect 6846 4326 6898 4378
rect 6910 4326 6962 4378
rect 4436 4224 4488 4276
rect 4896 4224 4948 4276
rect 3516 4156 3568 4208
rect 6092 4224 6144 4276
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 4160 4020 4212 4072
rect 4804 4088 4856 4140
rect 4528 4020 4580 4072
rect 5080 4020 5132 4072
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5816 4088 5868 4140
rect 6000 4088 6052 4140
rect 3700 3884 3752 3936
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 5632 3952 5684 4004
rect 6460 3952 6512 4004
rect 1663 3782 1715 3834
rect 1727 3782 1779 3834
rect 1791 3782 1843 3834
rect 1855 3782 1907 3834
rect 1919 3782 1971 3834
rect 3089 3782 3141 3834
rect 3153 3782 3205 3834
rect 3217 3782 3269 3834
rect 3281 3782 3333 3834
rect 3345 3782 3397 3834
rect 4515 3782 4567 3834
rect 4579 3782 4631 3834
rect 4643 3782 4695 3834
rect 4707 3782 4759 3834
rect 4771 3782 4823 3834
rect 5941 3782 5993 3834
rect 6005 3782 6057 3834
rect 6069 3782 6121 3834
rect 6133 3782 6185 3834
rect 6197 3782 6249 3834
rect 3976 3680 4028 3732
rect 4712 3680 4764 3732
rect 5632 3680 5684 3732
rect 5816 3680 5868 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 6276 3680 6328 3732
rect 4896 3612 4948 3664
rect 3884 3544 3936 3596
rect 940 3408 992 3460
rect 4436 3544 4488 3596
rect 5724 3612 5776 3664
rect 4160 3476 4212 3528
rect 4620 3476 4672 3528
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 5080 3476 5132 3528
rect 4160 3340 4212 3392
rect 4252 3340 4304 3392
rect 5356 3476 5408 3528
rect 5540 3476 5592 3528
rect 6092 3476 6144 3528
rect 2376 3238 2428 3290
rect 2440 3238 2492 3290
rect 2504 3238 2556 3290
rect 2568 3238 2620 3290
rect 2632 3238 2684 3290
rect 3802 3238 3854 3290
rect 3866 3238 3918 3290
rect 3930 3238 3982 3290
rect 3994 3238 4046 3290
rect 4058 3238 4110 3290
rect 5228 3238 5280 3290
rect 5292 3238 5344 3290
rect 5356 3238 5408 3290
rect 5420 3238 5472 3290
rect 5484 3238 5536 3290
rect 6654 3238 6706 3290
rect 6718 3238 6770 3290
rect 6782 3238 6834 3290
rect 6846 3238 6898 3290
rect 6910 3238 6962 3290
rect 2872 3136 2924 3188
rect 4528 3136 4580 3188
rect 4712 3136 4764 3188
rect 5632 3136 5684 3188
rect 5264 3068 5316 3120
rect 5356 3111 5408 3120
rect 5356 3077 5365 3111
rect 5365 3077 5399 3111
rect 5399 3077 5408 3111
rect 5356 3068 5408 3077
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 4804 2796 4856 2848
rect 4988 3000 5040 3052
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 6000 3068 6052 3120
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 5816 2864 5868 2916
rect 6368 2932 6420 2984
rect 1663 2694 1715 2746
rect 1727 2694 1779 2746
rect 1791 2694 1843 2746
rect 1855 2694 1907 2746
rect 1919 2694 1971 2746
rect 3089 2694 3141 2746
rect 3153 2694 3205 2746
rect 3217 2694 3269 2746
rect 3281 2694 3333 2746
rect 3345 2694 3397 2746
rect 4515 2694 4567 2746
rect 4579 2694 4631 2746
rect 4643 2694 4695 2746
rect 4707 2694 4759 2746
rect 4771 2694 4823 2746
rect 5941 2694 5993 2746
rect 6005 2694 6057 2746
rect 6069 2694 6121 2746
rect 6133 2694 6185 2746
rect 6197 2694 6249 2746
rect 5080 2592 5132 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 2780 2388 2832 2440
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6184 2456 6236 2508
rect 1584 2363 1636 2372
rect 1584 2329 1593 2363
rect 1593 2329 1627 2363
rect 1627 2329 1636 2363
rect 1584 2320 1636 2329
rect 5356 2320 5408 2372
rect 5080 2252 5132 2304
rect 2376 2150 2428 2202
rect 2440 2150 2492 2202
rect 2504 2150 2556 2202
rect 2568 2150 2620 2202
rect 2632 2150 2684 2202
rect 3802 2150 3854 2202
rect 3866 2150 3918 2202
rect 3930 2150 3982 2202
rect 3994 2150 4046 2202
rect 4058 2150 4110 2202
rect 5228 2150 5280 2202
rect 5292 2150 5344 2202
rect 5356 2150 5408 2202
rect 5420 2150 5472 2202
rect 5484 2150 5536 2202
rect 6654 2150 6706 2202
rect 6718 2150 6770 2202
rect 6782 2150 6834 2202
rect 6846 2150 6898 2202
rect 6910 2150 6962 2202
rect 4160 2048 4212 2100
rect 5816 2048 5868 2100
<< metal2 >>
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2376 5468 2684 5477
rect 2376 5466 2382 5468
rect 2438 5466 2462 5468
rect 2518 5466 2542 5468
rect 2598 5466 2622 5468
rect 2678 5466 2684 5468
rect 2438 5414 2440 5466
rect 2620 5414 2622 5466
rect 2376 5412 2382 5414
rect 2438 5412 2462 5414
rect 2518 5412 2542 5414
rect 2598 5412 2622 5414
rect 2678 5412 2684 5414
rect 2376 5403 2684 5412
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 940 5160 992 5166
rect 2700 5137 2728 5170
rect 940 5102 992 5108
rect 2686 5128 2742 5137
rect 952 5001 980 5102
rect 2686 5063 2742 5072
rect 938 4992 994 5001
rect 938 4927 994 4936
rect 1663 4924 1971 4933
rect 1663 4922 1669 4924
rect 1725 4922 1749 4924
rect 1805 4922 1829 4924
rect 1885 4922 1909 4924
rect 1965 4922 1971 4924
rect 1725 4870 1727 4922
rect 1907 4870 1909 4922
rect 1663 4868 1669 4870
rect 1725 4868 1749 4870
rect 1805 4868 1829 4870
rect 1885 4868 1909 4870
rect 1965 4868 1971 4870
rect 1663 4859 1971 4868
rect 2792 4690 2820 6831
rect 3514 6080 3570 6089
rect 3436 6038 3514 6066
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2596 4616 2648 4622
rect 2686 4584 2742 4593
rect 2648 4564 2686 4570
rect 2596 4558 2686 4564
rect 2608 4542 2686 4558
rect 2686 4519 2742 4528
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2376 4380 2684 4389
rect 2376 4378 2382 4380
rect 2438 4378 2462 4380
rect 2518 4378 2542 4380
rect 2598 4378 2622 4380
rect 2678 4378 2684 4380
rect 2438 4326 2440 4378
rect 2620 4326 2622 4378
rect 2376 4324 2382 4326
rect 2438 4324 2462 4326
rect 2518 4324 2542 4326
rect 2598 4324 2622 4326
rect 2678 4324 2684 4326
rect 2376 4315 2684 4324
rect 1663 3836 1971 3845
rect 1663 3834 1669 3836
rect 1725 3834 1749 3836
rect 1805 3834 1829 3836
rect 1885 3834 1909 3836
rect 1965 3834 1971 3836
rect 1725 3782 1727 3834
rect 1907 3782 1909 3834
rect 1663 3780 1669 3782
rect 1725 3780 1749 3782
rect 1805 3780 1829 3782
rect 1885 3780 1909 3782
rect 1965 3780 1971 3782
rect 1663 3771 1971 3780
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3097 980 3402
rect 2376 3292 2684 3301
rect 2376 3290 2382 3292
rect 2438 3290 2462 3292
rect 2518 3290 2542 3292
rect 2598 3290 2622 3292
rect 2678 3290 2684 3292
rect 2438 3238 2440 3290
rect 2620 3238 2622 3290
rect 2376 3236 2382 3238
rect 2438 3236 2462 3238
rect 2518 3236 2542 3238
rect 2598 3236 2622 3238
rect 2678 3236 2684 3238
rect 2376 3227 2684 3236
rect 938 3088 994 3097
rect 938 3023 994 3032
rect 1663 2748 1971 2757
rect 1663 2746 1669 2748
rect 1725 2746 1749 2748
rect 1805 2746 1829 2748
rect 1885 2746 1909 2748
rect 1965 2746 1971 2748
rect 1725 2694 1727 2746
rect 1907 2694 1909 2746
rect 1663 2692 1669 2694
rect 1725 2692 1749 2694
rect 1805 2692 1829 2694
rect 1885 2692 1909 2694
rect 1965 2692 1971 2694
rect 1663 2683 1971 2692
rect 2792 2446 2820 4490
rect 2884 3194 2912 5034
rect 2976 4690 3004 5850
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3344 5234 3372 5714
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3089 4924 3397 4933
rect 3089 4922 3095 4924
rect 3151 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3397 4924
rect 3151 4870 3153 4922
rect 3333 4870 3335 4922
rect 3089 4868 3095 4870
rect 3151 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3397 4870
rect 3089 4859 3397 4868
rect 3332 4752 3384 4758
rect 3330 4720 3332 4729
rect 3384 4720 3386 4729
rect 2964 4684 3016 4690
rect 3330 4655 3386 4664
rect 2964 4626 3016 4632
rect 3436 4622 3464 6038
rect 3514 6015 3570 6024
rect 6552 5840 6604 5846
rect 3514 5808 3570 5817
rect 6552 5782 6604 5788
rect 3514 5743 3570 5752
rect 3528 5370 3556 5743
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3514 5264 3570 5273
rect 3620 5234 3648 5578
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3514 5199 3516 5208
rect 3568 5199 3570 5208
rect 3608 5228 3660 5234
rect 3516 5170 3568 5176
rect 3608 5170 3660 5176
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3528 4214 3556 4966
rect 3608 4752 3660 4758
rect 3712 4706 3740 5510
rect 3802 5468 4110 5477
rect 3802 5466 3808 5468
rect 3864 5466 3888 5468
rect 3944 5466 3968 5468
rect 4024 5466 4048 5468
rect 4104 5466 4110 5468
rect 3864 5414 3866 5466
rect 4046 5414 4048 5466
rect 3802 5412 3808 5414
rect 3864 5412 3888 5414
rect 3944 5412 3968 5414
rect 4024 5412 4048 5414
rect 4104 5412 4110 5414
rect 3802 5403 4110 5412
rect 3792 5364 3844 5370
rect 4172 5352 4200 5646
rect 5228 5468 5536 5477
rect 5228 5466 5234 5468
rect 5290 5466 5314 5468
rect 5370 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5536 5468
rect 5290 5414 5292 5466
rect 5472 5414 5474 5466
rect 5228 5412 5234 5414
rect 5290 5412 5314 5414
rect 5370 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5536 5414
rect 5228 5403 5536 5412
rect 3792 5306 3844 5312
rect 3988 5324 4200 5352
rect 4344 5364 4396 5370
rect 3804 5001 3832 5306
rect 3988 5234 4016 5324
rect 4344 5306 4396 5312
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 3976 5228 4028 5234
rect 4356 5216 4384 5306
rect 3976 5170 4028 5176
rect 4172 5188 4384 5216
rect 3790 4992 3846 5001
rect 3790 4927 3846 4936
rect 3988 4826 4016 5170
rect 4172 5114 4200 5188
rect 4080 5086 4200 5114
rect 4344 5092 4396 5098
rect 4080 4826 4108 5086
rect 4344 5034 4396 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4172 4826 4200 4966
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3660 4700 3740 4706
rect 3608 4694 3740 4700
rect 3620 4678 3740 4694
rect 3712 4622 3740 4678
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3712 3942 3740 4558
rect 3802 4380 4110 4389
rect 3802 4378 3808 4380
rect 3864 4378 3888 4380
rect 3944 4378 3968 4380
rect 4024 4378 4048 4380
rect 4104 4378 4110 4380
rect 3864 4326 3866 4378
rect 4046 4326 4048 4378
rect 3802 4324 3808 4326
rect 3864 4324 3888 4326
rect 3944 4324 3968 4326
rect 4024 4324 4048 4326
rect 4104 4324 4110 4326
rect 3802 4315 4110 4324
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3089 3836 3397 3845
rect 3089 3834 3095 3836
rect 3151 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3397 3836
rect 3151 3782 3153 3834
rect 3333 3782 3335 3834
rect 3089 3780 3095 3782
rect 3151 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3397 3782
rect 3089 3771 3397 3780
rect 3896 3602 3924 3878
rect 3988 3738 4016 3878
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 4080 3482 4108 4111
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4172 3641 4200 4014
rect 4158 3632 4214 3641
rect 4158 3567 4214 3576
rect 4160 3528 4212 3534
rect 4080 3476 4160 3482
rect 4080 3470 4212 3476
rect 4080 3454 4200 3470
rect 4264 3398 4292 4966
rect 4356 4622 4384 5034
rect 4448 4622 4476 5306
rect 5172 5296 5224 5302
rect 5000 5244 5172 5250
rect 5000 5238 5224 5244
rect 5000 5234 5212 5238
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4988 5228 5212 5234
rect 5040 5222 5212 5228
rect 4988 5170 5040 5176
rect 4540 5098 4568 5170
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4515 4924 4823 4933
rect 4515 4922 4521 4924
rect 4577 4922 4601 4924
rect 4657 4922 4681 4924
rect 4737 4922 4761 4924
rect 4817 4922 4823 4924
rect 4577 4870 4579 4922
rect 4759 4870 4761 4922
rect 4515 4868 4521 4870
rect 4577 4868 4601 4870
rect 4657 4868 4681 4870
rect 4737 4868 4761 4870
rect 4817 4868 4823 4870
rect 4515 4859 4823 4868
rect 4712 4820 4764 4826
rect 4908 4808 4936 5034
rect 4988 5024 5040 5030
rect 4986 4992 4988 5001
rect 5040 4992 5042 5001
rect 4986 4927 5042 4936
rect 5092 4808 5120 5102
rect 5184 4826 5212 5222
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 4712 4762 4764 4768
rect 4816 4780 4936 4808
rect 5000 4780 5120 4808
rect 5172 4820 5224 4826
rect 4724 4622 4752 4762
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4342 4448 4398 4457
rect 4342 4383 4398 4392
rect 4356 4146 4384 4383
rect 4448 4282 4476 4558
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4540 4078 4568 4422
rect 4528 4072 4580 4078
rect 4632 4049 4660 4422
rect 4816 4321 4844 4780
rect 5000 4570 5028 4780
rect 5172 4762 5224 4768
rect 5276 4672 5304 5170
rect 5368 4826 5396 5170
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5460 4758 5488 4966
rect 5552 4865 5580 5170
rect 5538 4856 5594 4865
rect 5538 4791 5594 4800
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 4908 4542 5028 4570
rect 5092 4644 5304 4672
rect 5540 4684 5592 4690
rect 4802 4312 4858 4321
rect 4908 4282 4936 4542
rect 4802 4247 4858 4256
rect 4896 4276 4948 4282
rect 4816 4146 4844 4247
rect 4896 4218 4948 4224
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 5092 4078 5120 4644
rect 5644 4672 5672 5646
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 5736 5234 5764 5510
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5920 5234 5948 5306
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5722 5128 5778 5137
rect 5722 5063 5778 5072
rect 5736 4826 5764 5063
rect 6276 5024 6328 5030
rect 6380 5001 6408 5510
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6276 4966 6328 4972
rect 6366 4992 6422 5001
rect 5941 4924 6249 4933
rect 5941 4922 5947 4924
rect 6003 4922 6027 4924
rect 6083 4922 6107 4924
rect 6163 4922 6187 4924
rect 6243 4922 6249 4924
rect 6003 4870 6005 4922
rect 6185 4870 6187 4922
rect 5941 4868 5947 4870
rect 6003 4868 6027 4870
rect 6083 4868 6107 4870
rect 6163 4868 6187 4870
rect 6243 4868 6249 4870
rect 5941 4859 6249 4868
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5592 4644 5672 4672
rect 5540 4626 5592 4632
rect 5170 4584 5226 4593
rect 5170 4519 5226 4528
rect 5184 4486 5212 4519
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5228 4380 5536 4389
rect 5228 4378 5234 4380
rect 5290 4378 5314 4380
rect 5370 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5536 4380
rect 5290 4326 5292 4378
rect 5472 4326 5474 4378
rect 5228 4324 5234 4326
rect 5290 4324 5314 4326
rect 5370 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5536 4326
rect 5228 4315 5536 4324
rect 5644 4146 5672 4644
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5080 4072 5132 4078
rect 4528 4014 4580 4020
rect 4618 4040 4674 4049
rect 5080 4014 5132 4020
rect 4618 3975 4674 3984
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 4515 3836 4823 3845
rect 4515 3834 4521 3836
rect 4577 3834 4601 3836
rect 4657 3834 4681 3836
rect 4737 3834 4761 3836
rect 4817 3834 4823 3836
rect 4577 3782 4579 3834
rect 4759 3782 4761 3834
rect 4515 3780 4521 3782
rect 4577 3780 4601 3782
rect 4657 3780 4681 3782
rect 4737 3780 4761 3782
rect 4817 3780 4823 3782
rect 4515 3771 4823 3780
rect 5644 3738 5672 3946
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 4436 3596 4488 3602
rect 4488 3556 4568 3584
rect 4436 3538 4488 3544
rect 4540 3505 4568 3556
rect 4620 3528 4672 3534
rect 4526 3496 4582 3505
rect 4620 3470 4672 3476
rect 4526 3431 4582 3440
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 3802 3292 4110 3301
rect 3802 3290 3808 3292
rect 3864 3290 3888 3292
rect 3944 3290 3968 3292
rect 4024 3290 4048 3292
rect 4104 3290 4110 3292
rect 3864 3238 3866 3290
rect 4046 3238 4048 3290
rect 3802 3236 3808 3238
rect 3864 3236 3888 3238
rect 3944 3236 3968 3238
rect 4024 3236 4048 3238
rect 4104 3236 4110 3238
rect 3802 3227 4110 3236
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3089 2748 3397 2757
rect 3089 2746 3095 2748
rect 3151 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3397 2748
rect 3151 2694 3153 2746
rect 3333 2694 3335 2746
rect 3089 2692 3095 2694
rect 3151 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3397 2694
rect 3089 2683 3397 2692
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1596 1329 1624 2314
rect 2376 2204 2684 2213
rect 2376 2202 2382 2204
rect 2438 2202 2462 2204
rect 2518 2202 2542 2204
rect 2598 2202 2622 2204
rect 2678 2202 2684 2204
rect 2438 2150 2440 2202
rect 2620 2150 2622 2202
rect 2376 2148 2382 2150
rect 2438 2148 2462 2150
rect 2518 2148 2542 2150
rect 2598 2148 2622 2150
rect 2678 2148 2684 2150
rect 2376 2139 2684 2148
rect 3802 2204 4110 2213
rect 3802 2202 3808 2204
rect 3864 2202 3888 2204
rect 3944 2202 3968 2204
rect 4024 2202 4048 2204
rect 4104 2202 4110 2204
rect 3864 2150 3866 2202
rect 4046 2150 4048 2202
rect 3802 2148 3808 2150
rect 3864 2148 3888 2150
rect 3944 2148 3968 2150
rect 4024 2148 4048 2150
rect 4104 2148 4110 2150
rect 3802 2139 4110 2148
rect 4172 2106 4200 3334
rect 4528 3188 4580 3194
rect 4632 3176 4660 3470
rect 4724 3194 4752 3674
rect 5736 3670 5764 4558
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5828 3738 5856 4082
rect 5920 4026 5948 4558
rect 6012 4146 6040 4694
rect 6288 4622 6316 4966
rect 6366 4927 6422 4936
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6104 4282 6132 4558
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5920 3998 6316 4026
rect 6472 4010 6500 5034
rect 6564 4729 6592 5782
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6654 5468 6962 5477
rect 6654 5466 6660 5468
rect 6716 5466 6740 5468
rect 6796 5466 6820 5468
rect 6876 5466 6900 5468
rect 6956 5466 6962 5468
rect 6716 5414 6718 5466
rect 6898 5414 6900 5466
rect 6654 5412 6660 5414
rect 6716 5412 6740 5414
rect 6796 5412 6820 5414
rect 6876 5412 6900 5414
rect 6956 5412 6962 5414
rect 6654 5403 6962 5412
rect 7024 5273 7052 5646
rect 7010 5264 7066 5273
rect 7010 5199 7066 5208
rect 6550 4720 6606 4729
rect 6550 4655 6606 4664
rect 6654 4380 6962 4389
rect 6654 4378 6660 4380
rect 6716 4378 6740 4380
rect 6796 4378 6820 4380
rect 6876 4378 6900 4380
rect 6956 4378 6962 4380
rect 6716 4326 6718 4378
rect 6898 4326 6900 4378
rect 6654 4324 6660 4326
rect 6716 4324 6740 4326
rect 6796 4324 6820 4326
rect 6876 4324 6900 4326
rect 6956 4324 6962 4326
rect 6654 4315 6962 4324
rect 5941 3836 6249 3845
rect 5941 3834 5947 3836
rect 6003 3834 6027 3836
rect 6083 3834 6107 3836
rect 6163 3834 6187 3836
rect 6243 3834 6249 3836
rect 6003 3782 6005 3834
rect 6185 3782 6187 3834
rect 5941 3780 5947 3782
rect 6003 3780 6027 3782
rect 6083 3780 6107 3782
rect 6163 3780 6187 3782
rect 6243 3780 6249 3782
rect 5941 3771 6249 3780
rect 6288 3738 6316 3998
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6366 3904 6422 3913
rect 6366 3839 6422 3848
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4580 3148 4660 3176
rect 4712 3188 4764 3194
rect 4528 3130 4580 3136
rect 4712 3130 4764 3136
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4264 2774 4292 2994
rect 4816 2938 4844 3470
rect 4908 3097 4936 3606
rect 5080 3528 5132 3534
rect 5356 3528 5408 3534
rect 5132 3488 5356 3516
rect 5080 3470 5132 3476
rect 5356 3470 5408 3476
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5092 3380 5120 3470
rect 5000 3352 5120 3380
rect 5552 3380 5580 3470
rect 5552 3352 5672 3380
rect 4894 3088 4950 3097
rect 5000 3058 5028 3352
rect 5228 3292 5536 3301
rect 5228 3290 5234 3292
rect 5290 3290 5314 3292
rect 5370 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5536 3292
rect 5290 3238 5292 3290
rect 5472 3238 5474 3290
rect 5228 3236 5234 3238
rect 5290 3236 5314 3238
rect 5370 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5536 3238
rect 5228 3227 5536 3236
rect 5644 3194 5672 3352
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 6012 3126 6040 3674
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 4894 3023 4950 3032
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 4816 2910 5028 2938
rect 4804 2848 4856 2854
rect 4856 2825 4936 2836
rect 4856 2816 4950 2825
rect 4856 2808 4894 2816
rect 4804 2790 4856 2796
rect 4264 2746 4476 2774
rect 4448 2553 4476 2746
rect 4515 2748 4823 2757
rect 4894 2751 4950 2760
rect 4515 2746 4521 2748
rect 4577 2746 4601 2748
rect 4657 2746 4681 2748
rect 4737 2746 4761 2748
rect 4817 2746 4823 2748
rect 4577 2694 4579 2746
rect 4759 2694 4761 2746
rect 4515 2692 4521 2694
rect 4577 2692 4601 2694
rect 4657 2692 4681 2694
rect 4737 2692 4761 2694
rect 4817 2692 4823 2694
rect 4515 2683 4823 2692
rect 4434 2544 4490 2553
rect 4434 2479 4490 2488
rect 5000 2258 5028 2910
rect 5092 2650 5120 2994
rect 5170 2952 5226 2961
rect 5170 2887 5226 2896
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5184 2446 5212 2887
rect 5276 2446 5304 3062
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5368 2378 5396 3062
rect 6104 3058 6132 3470
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6380 2990 6408 3839
rect 6654 3292 6962 3301
rect 6654 3290 6660 3292
rect 6716 3290 6740 3292
rect 6796 3290 6820 3292
rect 6876 3290 6900 3292
rect 6956 3290 6962 3292
rect 6716 3238 6718 3290
rect 6898 3238 6900 3290
rect 6654 3236 6660 3238
rect 6716 3236 6740 3238
rect 6796 3236 6820 3238
rect 6876 3236 6900 3238
rect 6956 3236 6962 3238
rect 6654 3227 6962 3236
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5630 2816 5686 2825
rect 5630 2751 5686 2760
rect 5644 2650 5672 2751
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5448 2440 5500 2446
rect 5828 2394 5856 2858
rect 5941 2748 6249 2757
rect 5941 2746 5947 2748
rect 6003 2746 6027 2748
rect 6083 2746 6107 2748
rect 6163 2746 6187 2748
rect 6243 2746 6249 2748
rect 6003 2694 6005 2746
rect 6185 2694 6187 2746
rect 5941 2692 5947 2694
rect 6003 2692 6027 2694
rect 6083 2692 6107 2694
rect 6163 2692 6187 2694
rect 6243 2692 6249 2694
rect 5941 2683 6249 2692
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6196 2417 6224 2450
rect 5500 2388 5856 2394
rect 5448 2382 5856 2388
rect 5356 2372 5408 2378
rect 5460 2366 5856 2382
rect 5356 2314 5408 2320
rect 5080 2304 5132 2310
rect 5000 2252 5080 2258
rect 5000 2246 5132 2252
rect 5000 2230 5120 2246
rect 5228 2204 5536 2213
rect 5228 2202 5234 2204
rect 5290 2202 5314 2204
rect 5370 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5536 2204
rect 5290 2150 5292 2202
rect 5472 2150 5474 2202
rect 5228 2148 5234 2150
rect 5290 2148 5314 2150
rect 5370 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5536 2150
rect 5228 2139 5536 2148
rect 5828 2106 5856 2366
rect 6182 2408 6238 2417
rect 6182 2343 6238 2352
rect 6654 2204 6962 2213
rect 6654 2202 6660 2204
rect 6716 2202 6740 2204
rect 6796 2202 6820 2204
rect 6876 2202 6900 2204
rect 6956 2202 6962 2204
rect 6716 2150 6718 2202
rect 6898 2150 6900 2202
rect 6654 2148 6660 2150
rect 6716 2148 6740 2150
rect 6796 2148 6820 2150
rect 6876 2148 6900 2150
rect 6956 2148 6962 2150
rect 6654 2139 6962 2148
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 1582 1320 1638 1329
rect 1582 1255 1638 1264
<< via2 >>
rect 2778 6840 2834 6896
rect 2382 5466 2438 5468
rect 2462 5466 2518 5468
rect 2542 5466 2598 5468
rect 2622 5466 2678 5468
rect 2382 5414 2428 5466
rect 2428 5414 2438 5466
rect 2462 5414 2492 5466
rect 2492 5414 2504 5466
rect 2504 5414 2518 5466
rect 2542 5414 2556 5466
rect 2556 5414 2568 5466
rect 2568 5414 2598 5466
rect 2622 5414 2632 5466
rect 2632 5414 2678 5466
rect 2382 5412 2438 5414
rect 2462 5412 2518 5414
rect 2542 5412 2598 5414
rect 2622 5412 2678 5414
rect 2686 5072 2742 5128
rect 938 4936 994 4992
rect 1669 4922 1725 4924
rect 1749 4922 1805 4924
rect 1829 4922 1885 4924
rect 1909 4922 1965 4924
rect 1669 4870 1715 4922
rect 1715 4870 1725 4922
rect 1749 4870 1779 4922
rect 1779 4870 1791 4922
rect 1791 4870 1805 4922
rect 1829 4870 1843 4922
rect 1843 4870 1855 4922
rect 1855 4870 1885 4922
rect 1909 4870 1919 4922
rect 1919 4870 1965 4922
rect 1669 4868 1725 4870
rect 1749 4868 1805 4870
rect 1829 4868 1885 4870
rect 1909 4868 1965 4870
rect 2686 4528 2742 4584
rect 2382 4378 2438 4380
rect 2462 4378 2518 4380
rect 2542 4378 2598 4380
rect 2622 4378 2678 4380
rect 2382 4326 2428 4378
rect 2428 4326 2438 4378
rect 2462 4326 2492 4378
rect 2492 4326 2504 4378
rect 2504 4326 2518 4378
rect 2542 4326 2556 4378
rect 2556 4326 2568 4378
rect 2568 4326 2598 4378
rect 2622 4326 2632 4378
rect 2632 4326 2678 4378
rect 2382 4324 2438 4326
rect 2462 4324 2518 4326
rect 2542 4324 2598 4326
rect 2622 4324 2678 4326
rect 1669 3834 1725 3836
rect 1749 3834 1805 3836
rect 1829 3834 1885 3836
rect 1909 3834 1965 3836
rect 1669 3782 1715 3834
rect 1715 3782 1725 3834
rect 1749 3782 1779 3834
rect 1779 3782 1791 3834
rect 1791 3782 1805 3834
rect 1829 3782 1843 3834
rect 1843 3782 1855 3834
rect 1855 3782 1885 3834
rect 1909 3782 1919 3834
rect 1919 3782 1965 3834
rect 1669 3780 1725 3782
rect 1749 3780 1805 3782
rect 1829 3780 1885 3782
rect 1909 3780 1965 3782
rect 2382 3290 2438 3292
rect 2462 3290 2518 3292
rect 2542 3290 2598 3292
rect 2622 3290 2678 3292
rect 2382 3238 2428 3290
rect 2428 3238 2438 3290
rect 2462 3238 2492 3290
rect 2492 3238 2504 3290
rect 2504 3238 2518 3290
rect 2542 3238 2556 3290
rect 2556 3238 2568 3290
rect 2568 3238 2598 3290
rect 2622 3238 2632 3290
rect 2632 3238 2678 3290
rect 2382 3236 2438 3238
rect 2462 3236 2518 3238
rect 2542 3236 2598 3238
rect 2622 3236 2678 3238
rect 938 3032 994 3088
rect 1669 2746 1725 2748
rect 1749 2746 1805 2748
rect 1829 2746 1885 2748
rect 1909 2746 1965 2748
rect 1669 2694 1715 2746
rect 1715 2694 1725 2746
rect 1749 2694 1779 2746
rect 1779 2694 1791 2746
rect 1791 2694 1805 2746
rect 1829 2694 1843 2746
rect 1843 2694 1855 2746
rect 1855 2694 1885 2746
rect 1909 2694 1919 2746
rect 1919 2694 1965 2746
rect 1669 2692 1725 2694
rect 1749 2692 1805 2694
rect 1829 2692 1885 2694
rect 1909 2692 1965 2694
rect 3095 4922 3151 4924
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3095 4870 3141 4922
rect 3141 4870 3151 4922
rect 3175 4870 3205 4922
rect 3205 4870 3217 4922
rect 3217 4870 3231 4922
rect 3255 4870 3269 4922
rect 3269 4870 3281 4922
rect 3281 4870 3311 4922
rect 3335 4870 3345 4922
rect 3345 4870 3391 4922
rect 3095 4868 3151 4870
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3330 4700 3332 4720
rect 3332 4700 3384 4720
rect 3384 4700 3386 4720
rect 3330 4664 3386 4700
rect 3514 6024 3570 6080
rect 3514 5752 3570 5808
rect 3514 5228 3570 5264
rect 3514 5208 3516 5228
rect 3516 5208 3568 5228
rect 3568 5208 3570 5228
rect 3808 5466 3864 5468
rect 3888 5466 3944 5468
rect 3968 5466 4024 5468
rect 4048 5466 4104 5468
rect 3808 5414 3854 5466
rect 3854 5414 3864 5466
rect 3888 5414 3918 5466
rect 3918 5414 3930 5466
rect 3930 5414 3944 5466
rect 3968 5414 3982 5466
rect 3982 5414 3994 5466
rect 3994 5414 4024 5466
rect 4048 5414 4058 5466
rect 4058 5414 4104 5466
rect 3808 5412 3864 5414
rect 3888 5412 3944 5414
rect 3968 5412 4024 5414
rect 4048 5412 4104 5414
rect 5234 5466 5290 5468
rect 5314 5466 5370 5468
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5234 5414 5280 5466
rect 5280 5414 5290 5466
rect 5314 5414 5344 5466
rect 5344 5414 5356 5466
rect 5356 5414 5370 5466
rect 5394 5414 5408 5466
rect 5408 5414 5420 5466
rect 5420 5414 5450 5466
rect 5474 5414 5484 5466
rect 5484 5414 5530 5466
rect 5234 5412 5290 5414
rect 5314 5412 5370 5414
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 3790 4936 3846 4992
rect 3808 4378 3864 4380
rect 3888 4378 3944 4380
rect 3968 4378 4024 4380
rect 4048 4378 4104 4380
rect 3808 4326 3854 4378
rect 3854 4326 3864 4378
rect 3888 4326 3918 4378
rect 3918 4326 3930 4378
rect 3930 4326 3944 4378
rect 3968 4326 3982 4378
rect 3982 4326 3994 4378
rect 3994 4326 4024 4378
rect 4048 4326 4058 4378
rect 4058 4326 4104 4378
rect 3808 4324 3864 4326
rect 3888 4324 3944 4326
rect 3968 4324 4024 4326
rect 4048 4324 4104 4326
rect 4066 4120 4122 4176
rect 3095 3834 3151 3836
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3095 3782 3141 3834
rect 3141 3782 3151 3834
rect 3175 3782 3205 3834
rect 3205 3782 3217 3834
rect 3217 3782 3231 3834
rect 3255 3782 3269 3834
rect 3269 3782 3281 3834
rect 3281 3782 3311 3834
rect 3335 3782 3345 3834
rect 3345 3782 3391 3834
rect 3095 3780 3151 3782
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 4158 3576 4214 3632
rect 4521 4922 4577 4924
rect 4601 4922 4657 4924
rect 4681 4922 4737 4924
rect 4761 4922 4817 4924
rect 4521 4870 4567 4922
rect 4567 4870 4577 4922
rect 4601 4870 4631 4922
rect 4631 4870 4643 4922
rect 4643 4870 4657 4922
rect 4681 4870 4695 4922
rect 4695 4870 4707 4922
rect 4707 4870 4737 4922
rect 4761 4870 4771 4922
rect 4771 4870 4817 4922
rect 4521 4868 4577 4870
rect 4601 4868 4657 4870
rect 4681 4868 4737 4870
rect 4761 4868 4817 4870
rect 4986 4972 4988 4992
rect 4988 4972 5040 4992
rect 5040 4972 5042 4992
rect 4986 4936 5042 4972
rect 4342 4392 4398 4448
rect 5538 4800 5594 4856
rect 4802 4256 4858 4312
rect 5722 5072 5778 5128
rect 5947 4922 6003 4924
rect 6027 4922 6083 4924
rect 6107 4922 6163 4924
rect 6187 4922 6243 4924
rect 5947 4870 5993 4922
rect 5993 4870 6003 4922
rect 6027 4870 6057 4922
rect 6057 4870 6069 4922
rect 6069 4870 6083 4922
rect 6107 4870 6121 4922
rect 6121 4870 6133 4922
rect 6133 4870 6163 4922
rect 6187 4870 6197 4922
rect 6197 4870 6243 4922
rect 5947 4868 6003 4870
rect 6027 4868 6083 4870
rect 6107 4868 6163 4870
rect 6187 4868 6243 4870
rect 5170 4528 5226 4584
rect 5234 4378 5290 4380
rect 5314 4378 5370 4380
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5234 4326 5280 4378
rect 5280 4326 5290 4378
rect 5314 4326 5344 4378
rect 5344 4326 5356 4378
rect 5356 4326 5370 4378
rect 5394 4326 5408 4378
rect 5408 4326 5420 4378
rect 5420 4326 5450 4378
rect 5474 4326 5484 4378
rect 5484 4326 5530 4378
rect 5234 4324 5290 4326
rect 5314 4324 5370 4326
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 4618 3984 4674 4040
rect 4521 3834 4577 3836
rect 4601 3834 4657 3836
rect 4681 3834 4737 3836
rect 4761 3834 4817 3836
rect 4521 3782 4567 3834
rect 4567 3782 4577 3834
rect 4601 3782 4631 3834
rect 4631 3782 4643 3834
rect 4643 3782 4657 3834
rect 4681 3782 4695 3834
rect 4695 3782 4707 3834
rect 4707 3782 4737 3834
rect 4761 3782 4771 3834
rect 4771 3782 4817 3834
rect 4521 3780 4577 3782
rect 4601 3780 4657 3782
rect 4681 3780 4737 3782
rect 4761 3780 4817 3782
rect 4526 3440 4582 3496
rect 3808 3290 3864 3292
rect 3888 3290 3944 3292
rect 3968 3290 4024 3292
rect 4048 3290 4104 3292
rect 3808 3238 3854 3290
rect 3854 3238 3864 3290
rect 3888 3238 3918 3290
rect 3918 3238 3930 3290
rect 3930 3238 3944 3290
rect 3968 3238 3982 3290
rect 3982 3238 3994 3290
rect 3994 3238 4024 3290
rect 4048 3238 4058 3290
rect 4058 3238 4104 3290
rect 3808 3236 3864 3238
rect 3888 3236 3944 3238
rect 3968 3236 4024 3238
rect 4048 3236 4104 3238
rect 3095 2746 3151 2748
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3095 2694 3141 2746
rect 3141 2694 3151 2746
rect 3175 2694 3205 2746
rect 3205 2694 3217 2746
rect 3217 2694 3231 2746
rect 3255 2694 3269 2746
rect 3269 2694 3281 2746
rect 3281 2694 3311 2746
rect 3335 2694 3345 2746
rect 3345 2694 3391 2746
rect 3095 2692 3151 2694
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 2382 2202 2438 2204
rect 2462 2202 2518 2204
rect 2542 2202 2598 2204
rect 2622 2202 2678 2204
rect 2382 2150 2428 2202
rect 2428 2150 2438 2202
rect 2462 2150 2492 2202
rect 2492 2150 2504 2202
rect 2504 2150 2518 2202
rect 2542 2150 2556 2202
rect 2556 2150 2568 2202
rect 2568 2150 2598 2202
rect 2622 2150 2632 2202
rect 2632 2150 2678 2202
rect 2382 2148 2438 2150
rect 2462 2148 2518 2150
rect 2542 2148 2598 2150
rect 2622 2148 2678 2150
rect 3808 2202 3864 2204
rect 3888 2202 3944 2204
rect 3968 2202 4024 2204
rect 4048 2202 4104 2204
rect 3808 2150 3854 2202
rect 3854 2150 3864 2202
rect 3888 2150 3918 2202
rect 3918 2150 3930 2202
rect 3930 2150 3944 2202
rect 3968 2150 3982 2202
rect 3982 2150 3994 2202
rect 3994 2150 4024 2202
rect 4048 2150 4058 2202
rect 4058 2150 4104 2202
rect 3808 2148 3864 2150
rect 3888 2148 3944 2150
rect 3968 2148 4024 2150
rect 4048 2148 4104 2150
rect 6366 4936 6422 4992
rect 6660 5466 6716 5468
rect 6740 5466 6796 5468
rect 6820 5466 6876 5468
rect 6900 5466 6956 5468
rect 6660 5414 6706 5466
rect 6706 5414 6716 5466
rect 6740 5414 6770 5466
rect 6770 5414 6782 5466
rect 6782 5414 6796 5466
rect 6820 5414 6834 5466
rect 6834 5414 6846 5466
rect 6846 5414 6876 5466
rect 6900 5414 6910 5466
rect 6910 5414 6956 5466
rect 6660 5412 6716 5414
rect 6740 5412 6796 5414
rect 6820 5412 6876 5414
rect 6900 5412 6956 5414
rect 7010 5208 7066 5264
rect 6550 4664 6606 4720
rect 6660 4378 6716 4380
rect 6740 4378 6796 4380
rect 6820 4378 6876 4380
rect 6900 4378 6956 4380
rect 6660 4326 6706 4378
rect 6706 4326 6716 4378
rect 6740 4326 6770 4378
rect 6770 4326 6782 4378
rect 6782 4326 6796 4378
rect 6820 4326 6834 4378
rect 6834 4326 6846 4378
rect 6846 4326 6876 4378
rect 6900 4326 6910 4378
rect 6910 4326 6956 4378
rect 6660 4324 6716 4326
rect 6740 4324 6796 4326
rect 6820 4324 6876 4326
rect 6900 4324 6956 4326
rect 5947 3834 6003 3836
rect 6027 3834 6083 3836
rect 6107 3834 6163 3836
rect 6187 3834 6243 3836
rect 5947 3782 5993 3834
rect 5993 3782 6003 3834
rect 6027 3782 6057 3834
rect 6057 3782 6069 3834
rect 6069 3782 6083 3834
rect 6107 3782 6121 3834
rect 6121 3782 6133 3834
rect 6133 3782 6163 3834
rect 6187 3782 6197 3834
rect 6197 3782 6243 3834
rect 5947 3780 6003 3782
rect 6027 3780 6083 3782
rect 6107 3780 6163 3782
rect 6187 3780 6243 3782
rect 6366 3848 6422 3904
rect 4894 3032 4950 3088
rect 5234 3290 5290 3292
rect 5314 3290 5370 3292
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5234 3238 5280 3290
rect 5280 3238 5290 3290
rect 5314 3238 5344 3290
rect 5344 3238 5356 3290
rect 5356 3238 5370 3290
rect 5394 3238 5408 3290
rect 5408 3238 5420 3290
rect 5420 3238 5450 3290
rect 5474 3238 5484 3290
rect 5484 3238 5530 3290
rect 5234 3236 5290 3238
rect 5314 3236 5370 3238
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 4894 2760 4950 2816
rect 4521 2746 4577 2748
rect 4601 2746 4657 2748
rect 4681 2746 4737 2748
rect 4761 2746 4817 2748
rect 4521 2694 4567 2746
rect 4567 2694 4577 2746
rect 4601 2694 4631 2746
rect 4631 2694 4643 2746
rect 4643 2694 4657 2746
rect 4681 2694 4695 2746
rect 4695 2694 4707 2746
rect 4707 2694 4737 2746
rect 4761 2694 4771 2746
rect 4771 2694 4817 2746
rect 4521 2692 4577 2694
rect 4601 2692 4657 2694
rect 4681 2692 4737 2694
rect 4761 2692 4817 2694
rect 4434 2488 4490 2544
rect 5170 2896 5226 2952
rect 6660 3290 6716 3292
rect 6740 3290 6796 3292
rect 6820 3290 6876 3292
rect 6900 3290 6956 3292
rect 6660 3238 6706 3290
rect 6706 3238 6716 3290
rect 6740 3238 6770 3290
rect 6770 3238 6782 3290
rect 6782 3238 6796 3290
rect 6820 3238 6834 3290
rect 6834 3238 6846 3290
rect 6846 3238 6876 3290
rect 6900 3238 6910 3290
rect 6910 3238 6956 3290
rect 6660 3236 6716 3238
rect 6740 3236 6796 3238
rect 6820 3236 6876 3238
rect 6900 3236 6956 3238
rect 5630 2760 5686 2816
rect 5947 2746 6003 2748
rect 6027 2746 6083 2748
rect 6107 2746 6163 2748
rect 6187 2746 6243 2748
rect 5947 2694 5993 2746
rect 5993 2694 6003 2746
rect 6027 2694 6057 2746
rect 6057 2694 6069 2746
rect 6069 2694 6083 2746
rect 6107 2694 6121 2746
rect 6121 2694 6133 2746
rect 6133 2694 6163 2746
rect 6187 2694 6197 2746
rect 6197 2694 6243 2746
rect 5947 2692 6003 2694
rect 6027 2692 6083 2694
rect 6107 2692 6163 2694
rect 6187 2692 6243 2694
rect 5234 2202 5290 2204
rect 5314 2202 5370 2204
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5234 2150 5280 2202
rect 5280 2150 5290 2202
rect 5314 2150 5344 2202
rect 5344 2150 5356 2202
rect 5356 2150 5370 2202
rect 5394 2150 5408 2202
rect 5408 2150 5420 2202
rect 5420 2150 5450 2202
rect 5474 2150 5484 2202
rect 5484 2150 5530 2202
rect 5234 2148 5290 2150
rect 5314 2148 5370 2150
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 6182 2352 6238 2408
rect 6660 2202 6716 2204
rect 6740 2202 6796 2204
rect 6820 2202 6876 2204
rect 6900 2202 6956 2204
rect 6660 2150 6706 2202
rect 6706 2150 6716 2202
rect 6740 2150 6770 2202
rect 6770 2150 6782 2202
rect 6782 2150 6796 2202
rect 6820 2150 6834 2202
rect 6834 2150 6846 2202
rect 6846 2150 6876 2202
rect 6900 2150 6910 2202
rect 6910 2150 6956 2202
rect 6660 2148 6716 2150
rect 6740 2148 6796 2150
rect 6820 2148 6876 2150
rect 6900 2148 6956 2150
rect 1582 1264 1638 1320
<< metal3 >>
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 3509 6082 3575 6085
rect 7200 6082 8000 6112
rect 3509 6080 8000 6082
rect 3509 6024 3514 6080
rect 3570 6024 8000 6080
rect 3509 6022 8000 6024
rect 3509 6019 3575 6022
rect 7200 5992 8000 6022
rect 3509 5810 3575 5813
rect 7200 5810 8000 5840
rect 3509 5808 8000 5810
rect 3509 5752 3514 5808
rect 3570 5752 8000 5808
rect 3509 5750 8000 5752
rect 3509 5747 3575 5750
rect 7200 5720 8000 5750
rect 6502 5614 7114 5674
rect 2372 5472 2688 5473
rect 2372 5408 2378 5472
rect 2442 5408 2458 5472
rect 2522 5408 2538 5472
rect 2602 5408 2618 5472
rect 2682 5408 2688 5472
rect 2372 5407 2688 5408
rect 3798 5472 4114 5473
rect 3798 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4114 5472
rect 3798 5407 4114 5408
rect 5224 5472 5540 5473
rect 5224 5408 5230 5472
rect 5294 5408 5310 5472
rect 5374 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5540 5472
rect 5224 5407 5540 5408
rect 6502 5402 6562 5614
rect 7054 5538 7114 5614
rect 7200 5538 8000 5568
rect 7054 5478 8000 5538
rect 6650 5472 6966 5473
rect 6650 5408 6656 5472
rect 6720 5408 6736 5472
rect 6800 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6966 5472
rect 7200 5448 8000 5478
rect 6650 5407 6966 5408
rect 5766 5342 6562 5402
rect 3509 5266 3575 5269
rect 5766 5266 5826 5342
rect 3509 5264 5826 5266
rect 3509 5208 3514 5264
rect 3570 5208 5826 5264
rect 3509 5206 5826 5208
rect 7005 5266 7071 5269
rect 7200 5266 8000 5296
rect 7005 5264 8000 5266
rect 7005 5208 7010 5264
rect 7066 5208 8000 5264
rect 7005 5206 8000 5208
rect 3509 5203 3575 5206
rect 7005 5203 7071 5206
rect 7200 5176 8000 5206
rect 2681 5130 2747 5133
rect 5717 5130 5783 5133
rect 2681 5128 5783 5130
rect 2681 5072 2686 5128
rect 2742 5072 5722 5128
rect 5778 5072 5783 5128
rect 2681 5070 5783 5072
rect 2681 5067 2747 5070
rect 5717 5067 5783 5070
rect 0 4994 800 5024
rect 933 4994 999 4997
rect 0 4992 999 4994
rect 0 4936 938 4992
rect 994 4936 999 4992
rect 0 4934 999 4936
rect 0 4904 800 4934
rect 933 4931 999 4934
rect 3785 4994 3851 4997
rect 4981 4996 5047 4997
rect 4286 4994 4292 4996
rect 3785 4992 4292 4994
rect 3785 4936 3790 4992
rect 3846 4936 4292 4992
rect 3785 4934 4292 4936
rect 3785 4931 3851 4934
rect 4286 4932 4292 4934
rect 4356 4932 4362 4996
rect 4981 4992 5028 4996
rect 5092 4994 5098 4996
rect 6361 4994 6427 4997
rect 7200 4994 8000 5024
rect 4981 4936 4986 4992
rect 4981 4932 5028 4936
rect 5092 4934 5138 4994
rect 6361 4992 8000 4994
rect 6361 4936 6366 4992
rect 6422 4936 8000 4992
rect 6361 4934 8000 4936
rect 5092 4932 5098 4934
rect 4981 4931 5047 4932
rect 6361 4931 6427 4934
rect 1659 4928 1975 4929
rect 1659 4864 1665 4928
rect 1729 4864 1745 4928
rect 1809 4864 1825 4928
rect 1889 4864 1905 4928
rect 1969 4864 1975 4928
rect 1659 4863 1975 4864
rect 3085 4928 3401 4929
rect 3085 4864 3091 4928
rect 3155 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3401 4928
rect 3085 4863 3401 4864
rect 4511 4928 4827 4929
rect 4511 4864 4517 4928
rect 4581 4864 4597 4928
rect 4661 4864 4677 4928
rect 4741 4864 4757 4928
rect 4821 4864 4827 4928
rect 4511 4863 4827 4864
rect 5937 4928 6253 4929
rect 5937 4864 5943 4928
rect 6007 4864 6023 4928
rect 6087 4864 6103 4928
rect 6167 4864 6183 4928
rect 6247 4864 6253 4928
rect 7200 4904 8000 4934
rect 5937 4863 6253 4864
rect 5533 4858 5599 4861
rect 5758 4858 5764 4860
rect 5533 4856 5764 4858
rect 5533 4800 5538 4856
rect 5594 4800 5764 4856
rect 5533 4798 5764 4800
rect 5533 4795 5599 4798
rect 5758 4796 5764 4798
rect 5828 4796 5834 4860
rect 3325 4722 3391 4725
rect 6545 4722 6611 4725
rect 7200 4722 8000 4752
rect 3325 4720 5458 4722
rect 3325 4664 3330 4720
rect 3386 4664 5458 4720
rect 3325 4662 5458 4664
rect 3325 4659 3391 4662
rect 2681 4586 2747 4589
rect 5165 4586 5231 4589
rect 2681 4584 5231 4586
rect 2681 4528 2686 4584
rect 2742 4528 5170 4584
rect 5226 4528 5231 4584
rect 2681 4526 5231 4528
rect 5398 4586 5458 4662
rect 6545 4720 8000 4722
rect 6545 4664 6550 4720
rect 6606 4664 8000 4720
rect 6545 4662 8000 4664
rect 6545 4659 6611 4662
rect 7200 4632 8000 4662
rect 5398 4526 7114 4586
rect 2681 4523 2747 4526
rect 5165 4523 5231 4526
rect 4337 4450 4403 4453
rect 5022 4450 5028 4452
rect 4337 4448 5028 4450
rect 4337 4392 4342 4448
rect 4398 4392 5028 4448
rect 4337 4390 5028 4392
rect 4337 4387 4403 4390
rect 5022 4388 5028 4390
rect 5092 4388 5098 4452
rect 7054 4450 7114 4526
rect 7200 4450 8000 4480
rect 7054 4390 8000 4450
rect 2372 4384 2688 4385
rect 2372 4320 2378 4384
rect 2442 4320 2458 4384
rect 2522 4320 2538 4384
rect 2602 4320 2618 4384
rect 2682 4320 2688 4384
rect 2372 4319 2688 4320
rect 3798 4384 4114 4385
rect 3798 4320 3804 4384
rect 3868 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4114 4384
rect 3798 4319 4114 4320
rect 5224 4384 5540 4385
rect 5224 4320 5230 4384
rect 5294 4320 5310 4384
rect 5374 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5540 4384
rect 5224 4319 5540 4320
rect 6650 4384 6966 4385
rect 6650 4320 6656 4384
rect 6720 4320 6736 4384
rect 6800 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6966 4384
rect 7200 4360 8000 4390
rect 6650 4319 6966 4320
rect 4286 4252 4292 4316
rect 4356 4314 4362 4316
rect 4797 4314 4863 4317
rect 4356 4312 4863 4314
rect 4356 4256 4802 4312
rect 4858 4256 4863 4312
rect 4356 4254 4863 4256
rect 4356 4252 4362 4254
rect 4797 4251 4863 4254
rect 4061 4178 4127 4181
rect 7200 4178 8000 4208
rect 4061 4176 8000 4178
rect 4061 4120 4066 4176
rect 4122 4120 8000 4176
rect 4061 4118 8000 4120
rect 4061 4115 4127 4118
rect 7200 4088 8000 4118
rect 4613 4042 4679 4045
rect 5758 4042 5764 4044
rect 4613 4040 5764 4042
rect 4613 3984 4618 4040
rect 4674 3984 5764 4040
rect 4613 3982 5764 3984
rect 4613 3979 4679 3982
rect 5758 3980 5764 3982
rect 5828 3980 5834 4044
rect 6361 3906 6427 3909
rect 7200 3906 8000 3936
rect 6361 3904 8000 3906
rect 6361 3848 6366 3904
rect 6422 3848 8000 3904
rect 6361 3846 8000 3848
rect 6361 3843 6427 3846
rect 1659 3840 1975 3841
rect 1659 3776 1665 3840
rect 1729 3776 1745 3840
rect 1809 3776 1825 3840
rect 1889 3776 1905 3840
rect 1969 3776 1975 3840
rect 1659 3775 1975 3776
rect 3085 3840 3401 3841
rect 3085 3776 3091 3840
rect 3155 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3401 3840
rect 3085 3775 3401 3776
rect 4511 3840 4827 3841
rect 4511 3776 4517 3840
rect 4581 3776 4597 3840
rect 4661 3776 4677 3840
rect 4741 3776 4757 3840
rect 4821 3776 4827 3840
rect 4511 3775 4827 3776
rect 5937 3840 6253 3841
rect 5937 3776 5943 3840
rect 6007 3776 6023 3840
rect 6087 3776 6103 3840
rect 6167 3776 6183 3840
rect 6247 3776 6253 3840
rect 7200 3816 8000 3846
rect 5937 3775 6253 3776
rect 4153 3634 4219 3637
rect 7200 3634 8000 3664
rect 4153 3632 8000 3634
rect 4153 3576 4158 3632
rect 4214 3576 8000 3632
rect 4153 3574 8000 3576
rect 4153 3571 4219 3574
rect 7200 3544 8000 3574
rect 4521 3498 4587 3501
rect 4521 3496 7114 3498
rect 4521 3440 4526 3496
rect 4582 3440 7114 3496
rect 4521 3438 7114 3440
rect 4521 3435 4587 3438
rect 7054 3362 7114 3438
rect 7200 3362 8000 3392
rect 7054 3302 8000 3362
rect 2372 3296 2688 3297
rect 2372 3232 2378 3296
rect 2442 3232 2458 3296
rect 2522 3232 2538 3296
rect 2602 3232 2618 3296
rect 2682 3232 2688 3296
rect 2372 3231 2688 3232
rect 3798 3296 4114 3297
rect 3798 3232 3804 3296
rect 3868 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4114 3296
rect 3798 3231 4114 3232
rect 5224 3296 5540 3297
rect 5224 3232 5230 3296
rect 5294 3232 5310 3296
rect 5374 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5540 3296
rect 5224 3231 5540 3232
rect 6650 3296 6966 3297
rect 6650 3232 6656 3296
rect 6720 3232 6736 3296
rect 6800 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6966 3296
rect 7200 3272 8000 3302
rect 6650 3231 6966 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 4889 3090 4955 3093
rect 7200 3090 8000 3120
rect 4889 3088 8000 3090
rect 4889 3032 4894 3088
rect 4950 3032 8000 3088
rect 4889 3030 8000 3032
rect 4889 3027 4955 3030
rect 7200 3000 8000 3030
rect 5165 2954 5231 2957
rect 5165 2952 6378 2954
rect 5165 2896 5170 2952
rect 5226 2896 6378 2952
rect 5165 2894 6378 2896
rect 5165 2891 5231 2894
rect 4889 2818 4955 2821
rect 5625 2818 5691 2821
rect 4889 2816 5691 2818
rect 4889 2760 4894 2816
rect 4950 2760 5630 2816
rect 5686 2760 5691 2816
rect 4889 2758 5691 2760
rect 6318 2818 6378 2894
rect 7200 2818 8000 2848
rect 6318 2758 8000 2818
rect 4889 2755 4955 2758
rect 5625 2755 5691 2758
rect 1659 2752 1975 2753
rect 1659 2688 1665 2752
rect 1729 2688 1745 2752
rect 1809 2688 1825 2752
rect 1889 2688 1905 2752
rect 1969 2688 1975 2752
rect 1659 2687 1975 2688
rect 3085 2752 3401 2753
rect 3085 2688 3091 2752
rect 3155 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3401 2752
rect 3085 2687 3401 2688
rect 4511 2752 4827 2753
rect 4511 2688 4517 2752
rect 4581 2688 4597 2752
rect 4661 2688 4677 2752
rect 4741 2688 4757 2752
rect 4821 2688 4827 2752
rect 4511 2687 4827 2688
rect 5937 2752 6253 2753
rect 5937 2688 5943 2752
rect 6007 2688 6023 2752
rect 6087 2688 6103 2752
rect 6167 2688 6183 2752
rect 6247 2688 6253 2752
rect 7200 2728 8000 2758
rect 5937 2687 6253 2688
rect 4429 2546 4495 2549
rect 7200 2546 8000 2576
rect 4429 2544 8000 2546
rect 4429 2488 4434 2544
rect 4490 2488 8000 2544
rect 4429 2486 8000 2488
rect 4429 2483 4495 2486
rect 7200 2456 8000 2486
rect 6177 2410 6243 2413
rect 6177 2408 7114 2410
rect 6177 2352 6182 2408
rect 6238 2352 7114 2408
rect 6177 2350 7114 2352
rect 6177 2347 6243 2350
rect 7054 2274 7114 2350
rect 7200 2274 8000 2304
rect 7054 2214 8000 2274
rect 2372 2208 2688 2209
rect 2372 2144 2378 2208
rect 2442 2144 2458 2208
rect 2522 2144 2538 2208
rect 2602 2144 2618 2208
rect 2682 2144 2688 2208
rect 2372 2143 2688 2144
rect 3798 2208 4114 2209
rect 3798 2144 3804 2208
rect 3868 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4114 2208
rect 3798 2143 4114 2144
rect 5224 2208 5540 2209
rect 5224 2144 5230 2208
rect 5294 2144 5310 2208
rect 5374 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5540 2208
rect 5224 2143 5540 2144
rect 6650 2208 6966 2209
rect 6650 2144 6656 2208
rect 6720 2144 6736 2208
rect 6800 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6966 2208
rect 7200 2184 8000 2214
rect 6650 2143 6966 2144
rect 7200 1912 8000 2032
rect 1577 1322 1643 1325
rect 798 1320 1643 1322
rect 798 1264 1582 1320
rect 1638 1264 1643 1320
rect 798 1262 1643 1264
rect 798 1216 858 1262
rect 1577 1259 1643 1262
rect 0 1126 858 1216
rect 0 1096 800 1126
<< via3 >>
rect 2378 5468 2442 5472
rect 2378 5412 2382 5468
rect 2382 5412 2438 5468
rect 2438 5412 2442 5468
rect 2378 5408 2442 5412
rect 2458 5468 2522 5472
rect 2458 5412 2462 5468
rect 2462 5412 2518 5468
rect 2518 5412 2522 5468
rect 2458 5408 2522 5412
rect 2538 5468 2602 5472
rect 2538 5412 2542 5468
rect 2542 5412 2598 5468
rect 2598 5412 2602 5468
rect 2538 5408 2602 5412
rect 2618 5468 2682 5472
rect 2618 5412 2622 5468
rect 2622 5412 2678 5468
rect 2678 5412 2682 5468
rect 2618 5408 2682 5412
rect 3804 5468 3868 5472
rect 3804 5412 3808 5468
rect 3808 5412 3864 5468
rect 3864 5412 3868 5468
rect 3804 5408 3868 5412
rect 3884 5468 3948 5472
rect 3884 5412 3888 5468
rect 3888 5412 3944 5468
rect 3944 5412 3948 5468
rect 3884 5408 3948 5412
rect 3964 5468 4028 5472
rect 3964 5412 3968 5468
rect 3968 5412 4024 5468
rect 4024 5412 4028 5468
rect 3964 5408 4028 5412
rect 4044 5468 4108 5472
rect 4044 5412 4048 5468
rect 4048 5412 4104 5468
rect 4104 5412 4108 5468
rect 4044 5408 4108 5412
rect 5230 5468 5294 5472
rect 5230 5412 5234 5468
rect 5234 5412 5290 5468
rect 5290 5412 5294 5468
rect 5230 5408 5294 5412
rect 5310 5468 5374 5472
rect 5310 5412 5314 5468
rect 5314 5412 5370 5468
rect 5370 5412 5374 5468
rect 5310 5408 5374 5412
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 6656 5468 6720 5472
rect 6656 5412 6660 5468
rect 6660 5412 6716 5468
rect 6716 5412 6720 5468
rect 6656 5408 6720 5412
rect 6736 5468 6800 5472
rect 6736 5412 6740 5468
rect 6740 5412 6796 5468
rect 6796 5412 6800 5468
rect 6736 5408 6800 5412
rect 6816 5468 6880 5472
rect 6816 5412 6820 5468
rect 6820 5412 6876 5468
rect 6876 5412 6880 5468
rect 6816 5408 6880 5412
rect 6896 5468 6960 5472
rect 6896 5412 6900 5468
rect 6900 5412 6956 5468
rect 6956 5412 6960 5468
rect 6896 5408 6960 5412
rect 4292 4932 4356 4996
rect 5028 4992 5092 4996
rect 5028 4936 5042 4992
rect 5042 4936 5092 4992
rect 5028 4932 5092 4936
rect 1665 4924 1729 4928
rect 1665 4868 1669 4924
rect 1669 4868 1725 4924
rect 1725 4868 1729 4924
rect 1665 4864 1729 4868
rect 1745 4924 1809 4928
rect 1745 4868 1749 4924
rect 1749 4868 1805 4924
rect 1805 4868 1809 4924
rect 1745 4864 1809 4868
rect 1825 4924 1889 4928
rect 1825 4868 1829 4924
rect 1829 4868 1885 4924
rect 1885 4868 1889 4924
rect 1825 4864 1889 4868
rect 1905 4924 1969 4928
rect 1905 4868 1909 4924
rect 1909 4868 1965 4924
rect 1965 4868 1969 4924
rect 1905 4864 1969 4868
rect 3091 4924 3155 4928
rect 3091 4868 3095 4924
rect 3095 4868 3151 4924
rect 3151 4868 3155 4924
rect 3091 4864 3155 4868
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 4517 4924 4581 4928
rect 4517 4868 4521 4924
rect 4521 4868 4577 4924
rect 4577 4868 4581 4924
rect 4517 4864 4581 4868
rect 4597 4924 4661 4928
rect 4597 4868 4601 4924
rect 4601 4868 4657 4924
rect 4657 4868 4661 4924
rect 4597 4864 4661 4868
rect 4677 4924 4741 4928
rect 4677 4868 4681 4924
rect 4681 4868 4737 4924
rect 4737 4868 4741 4924
rect 4677 4864 4741 4868
rect 4757 4924 4821 4928
rect 4757 4868 4761 4924
rect 4761 4868 4817 4924
rect 4817 4868 4821 4924
rect 4757 4864 4821 4868
rect 5943 4924 6007 4928
rect 5943 4868 5947 4924
rect 5947 4868 6003 4924
rect 6003 4868 6007 4924
rect 5943 4864 6007 4868
rect 6023 4924 6087 4928
rect 6023 4868 6027 4924
rect 6027 4868 6083 4924
rect 6083 4868 6087 4924
rect 6023 4864 6087 4868
rect 6103 4924 6167 4928
rect 6103 4868 6107 4924
rect 6107 4868 6163 4924
rect 6163 4868 6167 4924
rect 6103 4864 6167 4868
rect 6183 4924 6247 4928
rect 6183 4868 6187 4924
rect 6187 4868 6243 4924
rect 6243 4868 6247 4924
rect 6183 4864 6247 4868
rect 5764 4796 5828 4860
rect 5028 4388 5092 4452
rect 2378 4380 2442 4384
rect 2378 4324 2382 4380
rect 2382 4324 2438 4380
rect 2438 4324 2442 4380
rect 2378 4320 2442 4324
rect 2458 4380 2522 4384
rect 2458 4324 2462 4380
rect 2462 4324 2518 4380
rect 2518 4324 2522 4380
rect 2458 4320 2522 4324
rect 2538 4380 2602 4384
rect 2538 4324 2542 4380
rect 2542 4324 2598 4380
rect 2598 4324 2602 4380
rect 2538 4320 2602 4324
rect 2618 4380 2682 4384
rect 2618 4324 2622 4380
rect 2622 4324 2678 4380
rect 2678 4324 2682 4380
rect 2618 4320 2682 4324
rect 3804 4380 3868 4384
rect 3804 4324 3808 4380
rect 3808 4324 3864 4380
rect 3864 4324 3868 4380
rect 3804 4320 3868 4324
rect 3884 4380 3948 4384
rect 3884 4324 3888 4380
rect 3888 4324 3944 4380
rect 3944 4324 3948 4380
rect 3884 4320 3948 4324
rect 3964 4380 4028 4384
rect 3964 4324 3968 4380
rect 3968 4324 4024 4380
rect 4024 4324 4028 4380
rect 3964 4320 4028 4324
rect 4044 4380 4108 4384
rect 4044 4324 4048 4380
rect 4048 4324 4104 4380
rect 4104 4324 4108 4380
rect 4044 4320 4108 4324
rect 5230 4380 5294 4384
rect 5230 4324 5234 4380
rect 5234 4324 5290 4380
rect 5290 4324 5294 4380
rect 5230 4320 5294 4324
rect 5310 4380 5374 4384
rect 5310 4324 5314 4380
rect 5314 4324 5370 4380
rect 5370 4324 5374 4380
rect 5310 4320 5374 4324
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 6656 4380 6720 4384
rect 6656 4324 6660 4380
rect 6660 4324 6716 4380
rect 6716 4324 6720 4380
rect 6656 4320 6720 4324
rect 6736 4380 6800 4384
rect 6736 4324 6740 4380
rect 6740 4324 6796 4380
rect 6796 4324 6800 4380
rect 6736 4320 6800 4324
rect 6816 4380 6880 4384
rect 6816 4324 6820 4380
rect 6820 4324 6876 4380
rect 6876 4324 6880 4380
rect 6816 4320 6880 4324
rect 6896 4380 6960 4384
rect 6896 4324 6900 4380
rect 6900 4324 6956 4380
rect 6956 4324 6960 4380
rect 6896 4320 6960 4324
rect 4292 4252 4356 4316
rect 5764 3980 5828 4044
rect 1665 3836 1729 3840
rect 1665 3780 1669 3836
rect 1669 3780 1725 3836
rect 1725 3780 1729 3836
rect 1665 3776 1729 3780
rect 1745 3836 1809 3840
rect 1745 3780 1749 3836
rect 1749 3780 1805 3836
rect 1805 3780 1809 3836
rect 1745 3776 1809 3780
rect 1825 3836 1889 3840
rect 1825 3780 1829 3836
rect 1829 3780 1885 3836
rect 1885 3780 1889 3836
rect 1825 3776 1889 3780
rect 1905 3836 1969 3840
rect 1905 3780 1909 3836
rect 1909 3780 1965 3836
rect 1965 3780 1969 3836
rect 1905 3776 1969 3780
rect 3091 3836 3155 3840
rect 3091 3780 3095 3836
rect 3095 3780 3151 3836
rect 3151 3780 3155 3836
rect 3091 3776 3155 3780
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 4517 3836 4581 3840
rect 4517 3780 4521 3836
rect 4521 3780 4577 3836
rect 4577 3780 4581 3836
rect 4517 3776 4581 3780
rect 4597 3836 4661 3840
rect 4597 3780 4601 3836
rect 4601 3780 4657 3836
rect 4657 3780 4661 3836
rect 4597 3776 4661 3780
rect 4677 3836 4741 3840
rect 4677 3780 4681 3836
rect 4681 3780 4737 3836
rect 4737 3780 4741 3836
rect 4677 3776 4741 3780
rect 4757 3836 4821 3840
rect 4757 3780 4761 3836
rect 4761 3780 4817 3836
rect 4817 3780 4821 3836
rect 4757 3776 4821 3780
rect 5943 3836 6007 3840
rect 5943 3780 5947 3836
rect 5947 3780 6003 3836
rect 6003 3780 6007 3836
rect 5943 3776 6007 3780
rect 6023 3836 6087 3840
rect 6023 3780 6027 3836
rect 6027 3780 6083 3836
rect 6083 3780 6087 3836
rect 6023 3776 6087 3780
rect 6103 3836 6167 3840
rect 6103 3780 6107 3836
rect 6107 3780 6163 3836
rect 6163 3780 6167 3836
rect 6103 3776 6167 3780
rect 6183 3836 6247 3840
rect 6183 3780 6187 3836
rect 6187 3780 6243 3836
rect 6243 3780 6247 3836
rect 6183 3776 6247 3780
rect 2378 3292 2442 3296
rect 2378 3236 2382 3292
rect 2382 3236 2438 3292
rect 2438 3236 2442 3292
rect 2378 3232 2442 3236
rect 2458 3292 2522 3296
rect 2458 3236 2462 3292
rect 2462 3236 2518 3292
rect 2518 3236 2522 3292
rect 2458 3232 2522 3236
rect 2538 3292 2602 3296
rect 2538 3236 2542 3292
rect 2542 3236 2598 3292
rect 2598 3236 2602 3292
rect 2538 3232 2602 3236
rect 2618 3292 2682 3296
rect 2618 3236 2622 3292
rect 2622 3236 2678 3292
rect 2678 3236 2682 3292
rect 2618 3232 2682 3236
rect 3804 3292 3868 3296
rect 3804 3236 3808 3292
rect 3808 3236 3864 3292
rect 3864 3236 3868 3292
rect 3804 3232 3868 3236
rect 3884 3292 3948 3296
rect 3884 3236 3888 3292
rect 3888 3236 3944 3292
rect 3944 3236 3948 3292
rect 3884 3232 3948 3236
rect 3964 3292 4028 3296
rect 3964 3236 3968 3292
rect 3968 3236 4024 3292
rect 4024 3236 4028 3292
rect 3964 3232 4028 3236
rect 4044 3292 4108 3296
rect 4044 3236 4048 3292
rect 4048 3236 4104 3292
rect 4104 3236 4108 3292
rect 4044 3232 4108 3236
rect 5230 3292 5294 3296
rect 5230 3236 5234 3292
rect 5234 3236 5290 3292
rect 5290 3236 5294 3292
rect 5230 3232 5294 3236
rect 5310 3292 5374 3296
rect 5310 3236 5314 3292
rect 5314 3236 5370 3292
rect 5370 3236 5374 3292
rect 5310 3232 5374 3236
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 6656 3292 6720 3296
rect 6656 3236 6660 3292
rect 6660 3236 6716 3292
rect 6716 3236 6720 3292
rect 6656 3232 6720 3236
rect 6736 3292 6800 3296
rect 6736 3236 6740 3292
rect 6740 3236 6796 3292
rect 6796 3236 6800 3292
rect 6736 3232 6800 3236
rect 6816 3292 6880 3296
rect 6816 3236 6820 3292
rect 6820 3236 6876 3292
rect 6876 3236 6880 3292
rect 6816 3232 6880 3236
rect 6896 3292 6960 3296
rect 6896 3236 6900 3292
rect 6900 3236 6956 3292
rect 6956 3236 6960 3292
rect 6896 3232 6960 3236
rect 1665 2748 1729 2752
rect 1665 2692 1669 2748
rect 1669 2692 1725 2748
rect 1725 2692 1729 2748
rect 1665 2688 1729 2692
rect 1745 2748 1809 2752
rect 1745 2692 1749 2748
rect 1749 2692 1805 2748
rect 1805 2692 1809 2748
rect 1745 2688 1809 2692
rect 1825 2748 1889 2752
rect 1825 2692 1829 2748
rect 1829 2692 1885 2748
rect 1885 2692 1889 2748
rect 1825 2688 1889 2692
rect 1905 2748 1969 2752
rect 1905 2692 1909 2748
rect 1909 2692 1965 2748
rect 1965 2692 1969 2748
rect 1905 2688 1969 2692
rect 3091 2748 3155 2752
rect 3091 2692 3095 2748
rect 3095 2692 3151 2748
rect 3151 2692 3155 2748
rect 3091 2688 3155 2692
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 4517 2748 4581 2752
rect 4517 2692 4521 2748
rect 4521 2692 4577 2748
rect 4577 2692 4581 2748
rect 4517 2688 4581 2692
rect 4597 2748 4661 2752
rect 4597 2692 4601 2748
rect 4601 2692 4657 2748
rect 4657 2692 4661 2748
rect 4597 2688 4661 2692
rect 4677 2748 4741 2752
rect 4677 2692 4681 2748
rect 4681 2692 4737 2748
rect 4737 2692 4741 2748
rect 4677 2688 4741 2692
rect 4757 2748 4821 2752
rect 4757 2692 4761 2748
rect 4761 2692 4817 2748
rect 4817 2692 4821 2748
rect 4757 2688 4821 2692
rect 5943 2748 6007 2752
rect 5943 2692 5947 2748
rect 5947 2692 6003 2748
rect 6003 2692 6007 2748
rect 5943 2688 6007 2692
rect 6023 2748 6087 2752
rect 6023 2692 6027 2748
rect 6027 2692 6083 2748
rect 6083 2692 6087 2748
rect 6023 2688 6087 2692
rect 6103 2748 6167 2752
rect 6103 2692 6107 2748
rect 6107 2692 6163 2748
rect 6163 2692 6167 2748
rect 6103 2688 6167 2692
rect 6183 2748 6247 2752
rect 6183 2692 6187 2748
rect 6187 2692 6243 2748
rect 6243 2692 6247 2748
rect 6183 2688 6247 2692
rect 2378 2204 2442 2208
rect 2378 2148 2382 2204
rect 2382 2148 2438 2204
rect 2438 2148 2442 2204
rect 2378 2144 2442 2148
rect 2458 2204 2522 2208
rect 2458 2148 2462 2204
rect 2462 2148 2518 2204
rect 2518 2148 2522 2204
rect 2458 2144 2522 2148
rect 2538 2204 2602 2208
rect 2538 2148 2542 2204
rect 2542 2148 2598 2204
rect 2598 2148 2602 2204
rect 2538 2144 2602 2148
rect 2618 2204 2682 2208
rect 2618 2148 2622 2204
rect 2622 2148 2678 2204
rect 2678 2148 2682 2204
rect 2618 2144 2682 2148
rect 3804 2204 3868 2208
rect 3804 2148 3808 2204
rect 3808 2148 3864 2204
rect 3864 2148 3868 2204
rect 3804 2144 3868 2148
rect 3884 2204 3948 2208
rect 3884 2148 3888 2204
rect 3888 2148 3944 2204
rect 3944 2148 3948 2204
rect 3884 2144 3948 2148
rect 3964 2204 4028 2208
rect 3964 2148 3968 2204
rect 3968 2148 4024 2204
rect 4024 2148 4028 2204
rect 3964 2144 4028 2148
rect 4044 2204 4108 2208
rect 4044 2148 4048 2204
rect 4048 2148 4104 2204
rect 4104 2148 4108 2204
rect 4044 2144 4108 2148
rect 5230 2204 5294 2208
rect 5230 2148 5234 2204
rect 5234 2148 5290 2204
rect 5290 2148 5294 2204
rect 5230 2144 5294 2148
rect 5310 2204 5374 2208
rect 5310 2148 5314 2204
rect 5314 2148 5370 2204
rect 5370 2148 5374 2204
rect 5310 2144 5374 2148
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 6656 2204 6720 2208
rect 6656 2148 6660 2204
rect 6660 2148 6716 2204
rect 6716 2148 6720 2204
rect 6656 2144 6720 2148
rect 6736 2204 6800 2208
rect 6736 2148 6740 2204
rect 6740 2148 6796 2204
rect 6796 2148 6800 2204
rect 6736 2144 6800 2148
rect 6816 2204 6880 2208
rect 6816 2148 6820 2204
rect 6820 2148 6876 2204
rect 6876 2148 6880 2204
rect 6816 2144 6880 2148
rect 6896 2204 6960 2208
rect 6896 2148 6900 2204
rect 6900 2148 6956 2204
rect 6956 2148 6960 2204
rect 6896 2144 6960 2148
<< metal4 >>
rect 1657 4928 1977 5488
rect 1657 4864 1665 4928
rect 1729 4864 1745 4928
rect 1809 4864 1825 4928
rect 1889 4864 1905 4928
rect 1969 4864 1977 4928
rect 1657 3840 1977 4864
rect 1657 3776 1665 3840
rect 1729 3776 1745 3840
rect 1809 3776 1825 3840
rect 1889 3776 1905 3840
rect 1969 3776 1977 3840
rect 1657 2752 1977 3776
rect 1657 2688 1665 2752
rect 1729 2688 1745 2752
rect 1809 2688 1825 2752
rect 1889 2688 1905 2752
rect 1969 2688 1977 2752
rect 1657 2128 1977 2688
rect 2370 5472 2690 5488
rect 2370 5408 2378 5472
rect 2442 5408 2458 5472
rect 2522 5408 2538 5472
rect 2602 5408 2618 5472
rect 2682 5408 2690 5472
rect 2370 4384 2690 5408
rect 2370 4320 2378 4384
rect 2442 4320 2458 4384
rect 2522 4320 2538 4384
rect 2602 4320 2618 4384
rect 2682 4320 2690 4384
rect 2370 3296 2690 4320
rect 2370 3232 2378 3296
rect 2442 3232 2458 3296
rect 2522 3232 2538 3296
rect 2602 3232 2618 3296
rect 2682 3232 2690 3296
rect 2370 2208 2690 3232
rect 2370 2144 2378 2208
rect 2442 2144 2458 2208
rect 2522 2144 2538 2208
rect 2602 2144 2618 2208
rect 2682 2144 2690 2208
rect 2370 2128 2690 2144
rect 3083 4928 3403 5488
rect 3083 4864 3091 4928
rect 3155 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3403 4928
rect 3083 3840 3403 4864
rect 3083 3776 3091 3840
rect 3155 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3403 3840
rect 3083 2752 3403 3776
rect 3083 2688 3091 2752
rect 3155 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3403 2752
rect 3083 2128 3403 2688
rect 3796 5472 4116 5488
rect 3796 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4116 5472
rect 3796 4384 4116 5408
rect 4291 4996 4357 4997
rect 4291 4932 4292 4996
rect 4356 4932 4357 4996
rect 4291 4931 4357 4932
rect 3796 4320 3804 4384
rect 3868 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4116 4384
rect 3796 3296 4116 4320
rect 4294 4317 4354 4931
rect 4509 4928 4829 5488
rect 5222 5472 5542 5488
rect 5222 5408 5230 5472
rect 5294 5408 5310 5472
rect 5374 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5542 5472
rect 5027 4996 5093 4997
rect 5027 4932 5028 4996
rect 5092 4932 5093 4996
rect 5027 4931 5093 4932
rect 4509 4864 4517 4928
rect 4581 4864 4597 4928
rect 4661 4864 4677 4928
rect 4741 4864 4757 4928
rect 4821 4864 4829 4928
rect 4291 4316 4357 4317
rect 4291 4252 4292 4316
rect 4356 4252 4357 4316
rect 4291 4251 4357 4252
rect 3796 3232 3804 3296
rect 3868 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4116 3296
rect 3796 2208 4116 3232
rect 3796 2144 3804 2208
rect 3868 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4116 2208
rect 3796 2128 4116 2144
rect 4509 3840 4829 4864
rect 5030 4453 5090 4931
rect 5027 4452 5093 4453
rect 5027 4388 5028 4452
rect 5092 4388 5093 4452
rect 5027 4387 5093 4388
rect 4509 3776 4517 3840
rect 4581 3776 4597 3840
rect 4661 3776 4677 3840
rect 4741 3776 4757 3840
rect 4821 3776 4829 3840
rect 4509 2752 4829 3776
rect 4509 2688 4517 2752
rect 4581 2688 4597 2752
rect 4661 2688 4677 2752
rect 4741 2688 4757 2752
rect 4821 2688 4829 2752
rect 4509 2128 4829 2688
rect 5222 4384 5542 5408
rect 5935 4928 6255 5488
rect 5935 4864 5943 4928
rect 6007 4864 6023 4928
rect 6087 4864 6103 4928
rect 6167 4864 6183 4928
rect 6247 4864 6255 4928
rect 5763 4860 5829 4861
rect 5763 4796 5764 4860
rect 5828 4796 5829 4860
rect 5763 4795 5829 4796
rect 5222 4320 5230 4384
rect 5294 4320 5310 4384
rect 5374 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5542 4384
rect 5222 3296 5542 4320
rect 5766 4045 5826 4795
rect 5763 4044 5829 4045
rect 5763 3980 5764 4044
rect 5828 3980 5829 4044
rect 5763 3979 5829 3980
rect 5222 3232 5230 3296
rect 5294 3232 5310 3296
rect 5374 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5542 3296
rect 5222 2208 5542 3232
rect 5222 2144 5230 2208
rect 5294 2144 5310 2208
rect 5374 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5542 2208
rect 5222 2128 5542 2144
rect 5935 3840 6255 4864
rect 5935 3776 5943 3840
rect 6007 3776 6023 3840
rect 6087 3776 6103 3840
rect 6167 3776 6183 3840
rect 6247 3776 6255 3840
rect 5935 2752 6255 3776
rect 5935 2688 5943 2752
rect 6007 2688 6023 2752
rect 6087 2688 6103 2752
rect 6167 2688 6183 2752
rect 6247 2688 6255 2752
rect 5935 2128 6255 2688
rect 6648 5472 6968 5488
rect 6648 5408 6656 5472
rect 6720 5408 6736 5472
rect 6800 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6968 5472
rect 6648 4384 6968 5408
rect 6648 4320 6656 4384
rect 6720 4320 6736 4384
rect 6800 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6968 4384
rect 6648 3296 6968 4320
rect 6648 3232 6656 3296
rect 6720 3232 6736 3296
rect 6800 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6968 3296
rect 6648 2208 6968 3232
rect 6648 2144 6656 2208
rect 6720 2144 6736 2208
rect 6800 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6968 2208
rect 6648 2128 6968 2144
use sky130_fd_sc_hd__inv_2  _16_
timestamp 1733718626
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _17_
timestamp 1733718626
transform -1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _18_
timestamp 1733718626
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _19_
timestamp 1733718626
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _20_
timestamp 1733718626
transform -1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _21_
timestamp 1733718626
transform 1 0 4968 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _22_
timestamp 1733718626
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _23_
timestamp 1733718626
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _24_
timestamp 1733718626
transform 1 0 5704 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _25_
timestamp 1733718626
transform -1 0 6072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _26_
timestamp 1733718626
transform -1 0 5244 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _27_
timestamp 1733718626
transform 1 0 5060 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _28_
timestamp 1733718626
transform -1 0 4416 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _29_
timestamp 1733718626
transform -1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _30_
timestamp 1733718626
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _31_
timestamp 1733718626
transform -1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _32_
timestamp 1733718626
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _33_
timestamp 1733718626
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _34_
timestamp 1733718626
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _35_
timestamp 1733718626
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19
timestamp 1733718626
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1733718626
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1733718626
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_37
timestamp 1733718626
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1733718626
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1733718626
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1733718626
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1733718626
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 1733718626
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_33
timestamp 1733718626
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1733718626
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1733718626
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1733718626
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1733718626
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1733718626
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1733718626
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 1733718626
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1733718626
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1733718626
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_38
timestamp 1733718626
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_57
timestamp 1733718626
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1733718626
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1733718626
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1733718626
transform 1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1733718626
transform 1 0 3772 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1733718626
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1733718626
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1733718626
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1733718626
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1733718626
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1733718626
transform -1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1733718626
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1733718626
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1733718626
transform 1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1733718626
transform -1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1733718626
transform -1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1733718626
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output16
timestamp 1733718626
transform -1 0 2852 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output17
timestamp 1733718626
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output18
timestamp 1733718626
transform -1 0 2852 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output19
timestamp 1733718626
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1733718626
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1733718626
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1733718626
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1733718626
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1733718626
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1733718626
transform -1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1733718626
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1733718626
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1733718626
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1733718626
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1733718626
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1733718626
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12
timestamp 1733718626
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1733718626
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1733718626
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1733718626
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1733718626
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1733718626
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1733718626
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1733718626
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
<< labels >>
flabel metal4 s 6648 2128 6968 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5222 2128 5542 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3796 2128 4116 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2370 2128 2690 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5935 2128 6255 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4509 2128 4829 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3083 2128 3403 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1657 2128 1977 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 7200 1912 8000 2032 0 FreeSans 600 0 0 0 in0
port 3 nsew
flabel metal3 s 7200 2184 8000 2304 0 FreeSans 600 0 0 0 in1
port 4 nsew
flabel metal3 s 7200 4632 8000 4752 0 FreeSans 600 0 0 0 in10
port 5 nsew
flabel metal3 s 7200 4904 8000 5024 0 FreeSans 600 0 0 0 in11
port 6 nsew
flabel metal3 s 7200 5176 8000 5296 0 FreeSans 600 0 0 0 in12
port 7 nsew
flabel metal3 s 7200 5448 8000 5568 0 FreeSans 600 0 0 0 in13
port 8 nsew
flabel metal3 s 7200 5720 8000 5840 0 FreeSans 600 0 0 0 in14
port 9 nsew
flabel metal3 s 7200 5992 8000 6112 0 FreeSans 600 0 0 0 in15
port 10 nsew
flabel metal3 s 7200 2456 8000 2576 0 FreeSans 600 0 0 0 in2
port 11 nsew
flabel metal3 s 7200 2728 8000 2848 0 FreeSans 600 0 0 0 in3
port 12 nsew
flabel metal3 s 7200 3000 8000 3120 0 FreeSans 600 0 0 0 in4
port 13 nsew
flabel metal3 s 7200 3272 8000 3392 0 FreeSans 600 0 0 0 in5
port 14 nsew
flabel metal3 s 7200 3544 8000 3664 0 FreeSans 600 0 0 0 in6
port 15 nsew
flabel metal3 s 7200 3816 8000 3936 0 FreeSans 600 0 0 0 in7
port 16 nsew
flabel metal3 s 7200 4088 8000 4208 0 FreeSans 600 0 0 0 in8
port 17 nsew
flabel metal3 s 7200 4360 8000 4480 0 FreeSans 600 0 0 0 in9
port 18 nsew
flabel metal3 s 0 1096 800 1216 0 FreeSans 600 0 0 0 out0
port 19 nsew
flabel metal3 s 0 3000 800 3120 0 FreeSans 600 0 0 0 out1
port 20 nsew
flabel metal3 s 0 4904 800 5024 0 FreeSans 600 0 0 0 out2
port 21 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 out3
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 8000 8000
<< end >>
