magic
tech sky130B
timestamp 1729956472
<< metal1 >>
rect 7410 -2500 7510 -2090
rect 11780 -2500 11880 -2090
rect 7410 -2600 11880 -2500
rect 7410 -4110 7510 -2600
rect 11780 -4110 11880 -2600
<< metal2 >>
rect 7130 2560 7370 2660
rect 10900 2560 11740 2660
rect 7130 1090 7370 1190
rect 10900 1090 11740 1190
rect 7130 -590 7370 -490
rect 10900 -590 11740 -490
rect 7130 -2060 7370 -1960
rect 10900 -2060 11740 -1960
rect 7130 -3780 7370 -3680
rect 10900 -3780 11740 -3680
rect 7130 -5250 7370 -5150
rect 10900 -5250 11740 -5150
rect 7130 -6930 7370 -6830
rect 10900 -6930 11740 -6830
rect 7130 -8400 7370 -8300
rect 10900 -8400 11740 -8300
<< metal3 >>
rect 8170 3640 8270 3880
rect 8860 3640 8960 3880
rect 10680 3640 10780 3880
rect 11370 3640 11470 3880
rect 12540 3640 12640 3870
rect 13230 3640 13330 3870
rect 15050 3640 15150 3870
rect 15740 3640 15840 3870
rect 7840 -2850 7940 -2420
rect 8170 -2700 8270 -1570
rect 8530 -2850 8630 -2420
rect 8860 -2700 8960 -1570
rect 10350 -2850 10450 -2420
rect 10680 -2700 10780 -1570
rect 11040 -2850 11140 -2420
rect 11370 -2700 11470 -1570
rect 12210 -2850 12310 -2420
rect 12540 -2700 12640 -1570
rect 12900 -2850 13000 -2420
rect 13230 -2700 13330 -1570
rect 14720 -2850 14820 -2420
rect 15050 -2700 15150 -1570
rect 15410 -2850 15510 -2420
rect 15740 -2700 15840 -1570
rect 7840 -9000 7940 -8760
rect 8530 -9000 8630 -8760
rect 10350 -9000 10450 -8760
rect 11040 -9000 11140 -8760
rect 12210 -8990 12310 -8760
rect 12900 -8990 13000 -8760
rect 14720 -8990 14820 -8760
rect 15410 -8990 15510 -8760
use 4x4crossbar  x1
timestamp 1729956472
transform 1 0 7470 0 1 440
box -200 -2960 4005 3300
use 4x4crossbar  x2
timestamp 1729956472
transform 1 0 11840 0 1 440
box -200 -2960 4005 3300
use 4x4crossbar  x3
timestamp 1729956472
transform 1 0 11840 0 1 -5900
box -200 -2960 4005 3300
use 4x4crossbar  x4
timestamp 1729956472
transform 1 0 7470 0 1 -5900
box -200 -2960 4005 3300
<< labels >>
flabel metal3 7840 -9000 7940 -8900 0 FreeSans 128 0 0 0 SL1
port 8 nsew
flabel metal3 8530 -9000 8630 -8900 0 FreeSans 128 0 0 0 SL2
port 17 nsew
flabel metal3 11040 -9000 11140 -8900 0 FreeSans 128 0 0 0 SL4
port 19 nsew
flabel metal2 7130 -8400 7230 -8300 0 FreeSans 128 0 0 0 WL8
port 16 nsew
flabel metal2 7130 -6930 7230 -6830 0 FreeSans 128 0 0 0 WL7
port 15 nsew
flabel metal2 7130 -5250 7230 -5150 0 FreeSans 128 0 0 0 WL6
port 14 nsew
flabel metal2 7130 -3780 7230 -3680 0 FreeSans 128 0 0 0 WL5
port 13 nsew
flabel metal3 10350 -9000 10450 -8900 0 FreeSans 128 0 0 0 SL3
port 18 nsew
flabel metal3 12210 -8990 12310 -8890 0 FreeSans 128 0 0 0 SL5
port 21 nsew
flabel metal3 12900 -8990 13000 -8890 0 FreeSans 128 0 0 0 SL6
port 22 nsew
flabel metal3 14720 -8990 14820 -8890 0 FreeSans 128 0 0 0 SL7
port 23 nsew
flabel metal3 15410 -8990 15510 -8890 0 FreeSans 128 0 0 0 SL8
port 24 nsew
flabel metal1 7410 -2600 7510 -2500 0 FreeSans 128 0 0 0 VSS
port 25 nsew
flabel metal2 7130 -2060 7230 -1960 0 FreeSans 128 0 0 0 WL4
port 12 nsew
flabel metal2 7130 -590 7230 -490 0 FreeSans 128 0 0 0 WL3
port 11 nsew
flabel metal2 7130 1090 7230 1190 0 FreeSans 128 0 0 0 WL2
port 10 nsew
flabel metal2 7130 2560 7230 2660 0 FreeSans 128 0 0 0 WL1
port 9 nsew
flabel metal3 10680 3780 10780 3880 0 FreeSans 128 0 0 0 BL3
port 2 nsew
flabel metal3 11370 3780 11470 3880 0 FreeSans 128 0 0 0 BL4
port 3 nsew
flabel metal3 12540 3770 12640 3870 0 FreeSans 128 0 0 0 BL5
port 4 nsew
flabel metal3 13230 3770 13330 3870 0 FreeSans 128 0 0 0 BL6
port 5 nsew
flabel metal3 15050 3770 15150 3870 0 FreeSans 128 0 0 0 BL7
port 6 nsew
flabel metal3 15740 3770 15840 3870 0 FreeSans 128 0 0 0 BL8
port 7 nsew
flabel metal3 8170 3780 8270 3880 0 FreeSans 128 0 0 0 BL1
port 0 nsew
flabel metal3 8860 3780 8960 3880 0 FreeSans 128 0 0 0 BL2
port 1 nsew
<< end >>
