magic
tech sky130B
magscale 1 2
timestamp 1733072092
<< nwell >>
rect -574 -1780 3812 1200
<< mvnsubdiff >>
rect -508 1122 3746 1134
rect -508 1022 -334 1122
rect 3572 1022 3746 1122
rect -508 1010 3746 1022
rect -508 960 -384 1010
rect -508 -1540 -496 960
rect -396 -1540 -384 960
rect -508 -1590 -384 -1540
rect 3622 960 3746 1010
rect 3622 -1540 3634 960
rect 3734 -1540 3746 960
rect 3622 -1590 3746 -1540
rect -508 -1602 3746 -1590
rect -508 -1702 -334 -1602
rect 3572 -1702 3746 -1602
rect -508 -1714 3746 -1702
<< mvnsubdiffcont >>
rect -334 1022 3572 1122
rect -496 -1540 -396 960
rect 3634 -1540 3734 960
rect -334 -1702 3572 -1602
<< locali >>
rect -496 960 -396 1122
rect -496 -1702 -396 -1540
rect 3634 960 3734 1122
rect 3634 -1702 3734 -1540
<< viali >>
rect -396 1022 -334 1122
rect -334 1022 3572 1122
rect 3572 1022 3634 1122
rect -496 -1471 -396 891
rect 3634 -1471 3734 891
rect -396 -1702 -334 -1602
rect -334 -1702 3572 -1602
rect 3572 -1702 3634 -1602
<< metal1 >>
rect -502 1122 3740 1128
rect -502 1022 -396 1122
rect 3634 1022 3740 1122
rect -502 1016 3740 1022
rect -502 891 -390 1016
rect -1936 -1298 -1836 -1198
rect -1946 -1568 -1846 -1468
rect -502 -1471 -496 891
rect -396 -1471 -390 891
rect 210 716 220 1016
rect 730 770 782 1016
rect 706 670 806 770
rect 3018 716 3028 1016
rect 3628 891 3740 1016
rect -110 492 -58 502
rect -110 -684 -58 440
rect 170 492 222 502
rect -26 398 26 408
rect -26 336 26 346
rect -18 246 18 336
rect -18 -308 18 -246
rect 60 -330 112 -30
rect -18 -470 18 -408
rect -18 -1052 18 -962
rect -26 -1062 26 -1052
rect -26 -1124 26 -1114
rect 60 -1300 112 -382
rect 170 -684 222 440
rect 450 492 502 502
rect 254 398 306 408
rect 254 336 306 346
rect 262 246 298 336
rect 262 -308 298 -246
rect 340 -330 392 -30
rect 262 -470 298 -408
rect 340 -682 392 -382
rect 450 -684 502 440
rect 730 492 782 670
rect 534 398 586 408
rect 534 336 586 346
rect 542 246 578 336
rect 542 -308 578 -246
rect 620 -330 672 -30
rect 542 -470 578 -408
rect 620 -682 672 -382
rect 730 -684 782 440
rect 1010 492 1062 502
rect 814 398 866 408
rect 814 336 866 346
rect 822 246 858 336
rect 822 -308 858 -246
rect 900 -330 952 -30
rect 822 -470 858 -408
rect 900 -682 952 -382
rect 1010 -684 1062 440
rect 1290 492 1342 502
rect 1094 398 1146 408
rect 1094 336 1146 346
rect 1102 246 1138 336
rect 1102 -308 1138 -246
rect 1180 -330 1232 -30
rect 1102 -470 1138 -408
rect 1180 -682 1232 -382
rect 1290 -684 1342 440
rect 1570 492 1622 502
rect 1374 398 1426 408
rect 1374 336 1426 346
rect 1382 246 1418 336
rect 1382 -308 1418 -246
rect 1460 -330 1512 -30
rect 1382 -470 1418 -408
rect 1460 -682 1512 -382
rect 1570 -684 1622 440
rect 1850 492 1902 502
rect 1654 398 1706 408
rect 1654 336 1706 346
rect 1662 246 1698 336
rect 1662 -308 1698 -246
rect 1740 -330 1792 -30
rect 1662 -470 1698 -408
rect 1740 -682 1792 -382
rect 1850 -684 1902 440
rect 2130 492 2182 502
rect 1934 398 1986 408
rect 1934 336 1986 346
rect 1942 246 1978 336
rect 1942 -308 1978 -246
rect 2020 -330 2072 -30
rect 1942 -470 1978 -408
rect 2020 -682 2072 -382
rect 2130 -684 2182 440
rect 2410 492 2462 502
rect 2214 398 2266 408
rect 2214 336 2266 346
rect 2222 246 2258 336
rect 2222 -308 2258 -246
rect 2300 -330 2352 -30
rect 2222 -470 2258 -408
rect 2300 -682 2352 -382
rect 2410 -684 2462 440
rect 2690 492 2742 502
rect 2494 398 2546 408
rect 2494 336 2546 346
rect 2502 246 2538 336
rect 2502 -308 2538 -246
rect 2580 -330 2632 -30
rect 2502 -470 2538 -408
rect 2580 -682 2632 -382
rect 2690 -684 2742 440
rect 2970 492 3022 502
rect 2774 398 2826 408
rect 2774 336 2826 346
rect 2782 246 2818 336
rect 2782 -308 2818 -246
rect 2860 -330 2912 -30
rect 2782 -470 2818 -408
rect 2860 -682 2912 -382
rect 2970 -684 3022 440
rect 3228 282 3238 290
rect 3062 246 3238 282
rect 3228 238 3238 246
rect 3290 238 3300 290
rect 3062 -308 3098 -246
rect 3140 -330 3192 -30
rect 3062 -470 3098 -408
rect 262 -1052 298 -962
rect 542 -1052 578 -962
rect 822 -1052 858 -962
rect 1102 -1052 1138 -962
rect 254 -1062 306 -1052
rect 254 -1124 306 -1114
rect 534 -1062 586 -1052
rect 534 -1124 586 -1114
rect 814 -1062 866 -1052
rect 814 -1124 866 -1114
rect 1094 -1062 1146 -1052
rect 1094 -1124 1146 -1114
rect 1382 -1168 1418 -962
rect 1662 -1168 1698 -962
rect 1942 -1052 1978 -962
rect 2222 -1052 2258 -962
rect 2502 -1052 2538 -962
rect 2782 -1052 2818 -962
rect 3062 -1052 3098 -962
rect 1934 -1062 1986 -1052
rect 1934 -1124 1986 -1114
rect 2214 -1062 2266 -1052
rect 2214 -1124 2266 -1114
rect 2494 -1062 2546 -1052
rect 2494 -1124 2546 -1114
rect 2774 -1062 2826 -1052
rect 2774 -1124 2826 -1114
rect 3054 -1062 3106 -1052
rect 3054 -1124 3106 -1114
rect 1374 -1178 1426 -1168
rect 1374 -1240 1426 -1230
rect 1654 -1178 1706 -1168
rect 1654 -1240 1706 -1230
rect -502 -1596 -390 -1471
rect 66 -1472 102 -1300
rect 404 -1472 414 -1462
rect 66 -1508 414 -1472
rect 404 -1514 414 -1508
rect 466 -1472 476 -1462
rect 1662 -1472 1698 -1240
rect 3140 -1372 3192 -382
rect 2468 -1424 2478 -1372
rect 2530 -1424 3192 -1372
rect 466 -1508 1698 -1472
rect 3628 -1471 3634 891
rect 3734 -1471 3740 891
rect 466 -1514 476 -1508
rect 3628 -1596 3740 -1471
rect -502 -1602 3740 -1596
rect -502 -1702 -396 -1602
rect 3634 -1702 3740 -1602
rect -502 -1708 3740 -1702
rect -1942 -1838 -1842 -1738
rect 890 -1824 942 -1814
rect 890 -1886 942 -1876
rect 2774 -1824 2826 -1814
rect 2774 -1886 2826 -1876
rect 330 -1912 382 -1902
rect 330 -1974 382 -1964
rect 610 -1912 662 -1902
rect 610 -1974 662 -1964
rect 178 -2012 230 -2002
rect 178 -2074 230 -2064
rect 186 -2360 222 -2074
rect 254 -2112 306 -2102
rect 254 -2174 306 -2164
rect 262 -2228 298 -2174
rect 338 -2360 374 -1974
rect 458 -2012 510 -2002
rect 458 -2074 510 -2064
rect 466 -2360 502 -2074
rect 534 -2112 586 -2102
rect 534 -2174 586 -2164
rect 542 -2228 578 -2174
rect 618 -2360 654 -1974
rect 814 -2112 866 -2102
rect 814 -2174 866 -2164
rect 822 -2228 858 -2174
rect 262 -2798 298 -2738
rect 542 -2798 578 -2738
rect 746 -2822 782 -2640
rect 822 -2798 858 -2738
rect 898 -2744 936 -1886
rect 1450 -1912 1502 -1902
rect 1450 -1974 1502 -1964
rect 1730 -1912 1782 -1902
rect 1730 -1974 1782 -1964
rect 2570 -1912 2622 -1902
rect 2570 -1974 2622 -1964
rect 1298 -2012 1350 -2002
rect 1298 -2074 1350 -2064
rect 1094 -2112 1146 -2102
rect 1094 -2174 1146 -2164
rect 1102 -2228 1138 -2174
rect 1306 -2360 1342 -2074
rect 1374 -2112 1426 -2102
rect 1374 -2174 1426 -2164
rect 1382 -2228 1418 -2174
rect 1458 -2360 1494 -1974
rect 1578 -2012 1630 -2002
rect 1578 -2074 1630 -2064
rect 1586 -2360 1622 -2074
rect 1654 -2112 1706 -2102
rect 1654 -2174 1706 -2164
rect 1662 -2228 1698 -2174
rect 1738 -2360 1774 -1974
rect 2418 -2012 2470 -2002
rect 2418 -2074 2470 -2064
rect 1934 -2112 1986 -2102
rect 1934 -2174 1986 -2164
rect 2214 -2112 2266 -2102
rect 2214 -2174 2266 -2164
rect 1942 -2228 1978 -2174
rect 2222 -2228 2258 -2174
rect 2426 -2360 2462 -2074
rect 2494 -2112 2546 -2102
rect 2494 -2174 2546 -2164
rect 2502 -2228 2538 -2174
rect 2578 -2360 2614 -1974
rect 2698 -2012 2750 -2002
rect 2698 -2074 2750 -2064
rect 2706 -2360 2742 -2074
rect 2782 -2102 2818 -1886
rect 2850 -1912 2902 -1902
rect 2850 -1974 2902 -1964
rect 2774 -2112 2826 -2102
rect 2774 -2174 2826 -2164
rect 2782 -2228 2818 -2174
rect 2858 -2360 2894 -1974
rect 178 -2836 230 -2826
rect 178 -2898 230 -2888
rect 458 -2836 510 -2826
rect 458 -2898 510 -2888
rect 738 -2832 790 -2822
rect 738 -2894 790 -2884
rect 186 -3178 222 -2898
rect 330 -2936 382 -2926
rect 330 -2998 382 -2988
rect 262 -3082 298 -3022
rect 338 -3180 374 -2998
rect 466 -3180 502 -2898
rect 898 -2926 934 -2744
rect 1026 -2822 1062 -2640
rect 1102 -2798 1138 -2738
rect 1018 -2832 1070 -2822
rect 1018 -2894 1070 -2884
rect 1178 -2926 1214 -2640
rect 1382 -2798 1418 -2738
rect 1662 -2798 1698 -2738
rect 1866 -2822 1902 -2640
rect 1942 -2798 1978 -2738
rect 1298 -2836 1350 -2826
rect 1298 -2898 1350 -2888
rect 1578 -2836 1630 -2826
rect 1578 -2898 1630 -2888
rect 1858 -2832 1910 -2822
rect 1858 -2894 1910 -2884
rect 610 -2936 662 -2926
rect 610 -2998 662 -2988
rect 890 -2936 942 -2926
rect 890 -2998 942 -2988
rect 1170 -2936 1222 -2926
rect 1170 -2998 1222 -2988
rect 542 -3082 578 -3022
rect 618 -3180 654 -2998
rect 822 -3082 858 -3022
rect 1102 -3082 1138 -3022
rect 1306 -3180 1342 -2898
rect 1450 -2936 1502 -2926
rect 1450 -2998 1502 -2988
rect 1382 -3082 1418 -3022
rect 262 -3646 298 -3592
rect 542 -3646 578 -3592
rect 254 -3656 306 -3646
rect 254 -3718 306 -3708
rect 534 -3656 586 -3646
rect 534 -3718 586 -3708
rect 746 -3846 782 -3460
rect 822 -3646 858 -3592
rect 814 -3656 866 -3646
rect 814 -3718 866 -3708
rect 898 -3746 934 -3460
rect 890 -3756 942 -3746
rect 890 -3818 942 -3808
rect 1026 -3846 1062 -3460
rect 1102 -3646 1138 -3592
rect 1094 -3656 1146 -3646
rect 1094 -3718 1146 -3708
rect 1178 -3746 1214 -3460
rect 1382 -3646 1418 -3592
rect 1374 -3656 1426 -3646
rect 1374 -3718 1426 -3708
rect 1170 -3756 1222 -3746
rect 1170 -3818 1222 -3808
rect 738 -3856 790 -3846
rect 738 -3918 790 -3908
rect 1018 -3856 1070 -3846
rect 1018 -3918 1070 -3908
rect 1458 -4018 1494 -2998
rect 1382 -4052 1494 -4018
rect 1382 -4362 1418 -4052
rect 1586 -4080 1622 -2898
rect 2018 -2926 2054 -2640
rect 2146 -2822 2182 -2640
rect 2222 -2798 2258 -2738
rect 2138 -2832 2190 -2822
rect 2138 -2894 2190 -2884
rect 2298 -2926 2334 -2640
rect 2502 -2798 2538 -2738
rect 2782 -2798 2818 -2738
rect 2418 -2836 2470 -2826
rect 2418 -2898 2470 -2888
rect 2698 -2836 2750 -2826
rect 2698 -2898 2750 -2888
rect 1730 -2936 1782 -2926
rect 1730 -2998 1782 -2988
rect 2010 -2936 2062 -2926
rect 2010 -2998 2062 -2988
rect 2290 -2936 2342 -2926
rect 2290 -2998 2342 -2988
rect 1662 -3082 1698 -3022
rect 1738 -3180 1774 -2998
rect 1942 -3082 1978 -3022
rect 2222 -3082 2258 -3022
rect 2426 -3180 2462 -2898
rect 2570 -2936 2622 -2926
rect 2570 -2998 2622 -2988
rect 2502 -3082 2538 -3022
rect 2578 -3180 2614 -2998
rect 2706 -3180 2742 -2898
rect 2850 -2936 2902 -2926
rect 2850 -2998 2902 -2988
rect 2782 -3082 2818 -3022
rect 2858 -3180 2894 -2998
rect 1662 -3646 1698 -3592
rect 1654 -3656 1706 -3646
rect 1654 -3718 1706 -3708
rect 1866 -3846 1902 -3460
rect 1942 -3646 1978 -3592
rect 1934 -3656 1986 -3646
rect 1934 -3718 1986 -3708
rect 2018 -3746 2054 -3460
rect 2010 -3756 2062 -3746
rect 2010 -3818 2062 -3808
rect 1858 -3856 1910 -3846
rect 1858 -3918 1910 -3908
rect 2018 -3946 2054 -3818
rect 2146 -3846 2182 -3460
rect 2222 -3646 2258 -3592
rect 2214 -3656 2266 -3646
rect 2214 -3718 2266 -3708
rect 2298 -3746 2334 -3460
rect 2502 -3646 2538 -3592
rect 2782 -3646 2818 -3592
rect 2494 -3656 2546 -3646
rect 2494 -3718 2546 -3708
rect 2774 -3656 2826 -3646
rect 2774 -3718 2826 -3708
rect 2290 -3756 2342 -3746
rect 2290 -3818 2342 -3808
rect 2138 -3856 2190 -3846
rect 2138 -3918 2190 -3908
rect 1458 -4116 1622 -4080
rect 1662 -3984 2054 -3946
rect 1458 -4118 1510 -4116
rect 1458 -4180 1510 -4170
rect 1458 -4450 1494 -4180
rect 1578 -4210 1630 -4200
rect 1578 -4272 1630 -4262
rect 1460 -4492 1494 -4450
rect 1584 -4494 1620 -4272
rect 1662 -4362 1698 -3984
rect 2148 -4028 2182 -3918
rect 1740 -4066 2182 -4028
rect 1304 -5028 1340 -4758
rect 1382 -4924 1418 -4838
rect 1480 -4872 1698 -4838
rect 1374 -4934 1426 -4924
rect 1374 -4996 1426 -4986
rect 1296 -5038 1348 -5028
rect 1480 -5032 1514 -4872
rect 1654 -4934 1706 -4924
rect 1654 -4996 1706 -4986
rect 1296 -5100 1348 -5090
rect 1382 -5066 1514 -5032
rect 1382 -5184 1418 -5066
rect 1458 -5118 1510 -5108
rect 1458 -5180 1510 -5170
rect 1458 -5296 1494 -5180
rect 1662 -5182 1698 -4996
rect 1740 -5014 1776 -4066
rect 1820 -4118 1872 -4108
rect 1820 -4180 1872 -4170
rect 1734 -5024 1786 -5014
rect 1734 -5086 1786 -5076
rect 1338 -5814 1374 -5642
rect 1584 -5718 1620 -5482
rect 1706 -5694 1742 -5482
rect 1822 -5694 1872 -4180
rect 1576 -5728 1628 -5718
rect 1706 -5730 1872 -5694
rect 1576 -5790 1628 -5780
rect 1330 -5824 1382 -5814
rect 1330 -5886 1382 -5876
rect 1338 -6014 1374 -5886
rect 1584 -6014 1620 -5790
<< via1 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -110 440 -58 492
rect 170 440 222 492
rect -26 346 26 398
rect 60 -382 112 -330
rect -26 -1114 26 -1062
rect 450 440 502 492
rect 254 346 306 398
rect 340 -382 392 -330
rect 730 440 782 492
rect 534 346 586 398
rect 620 -382 672 -330
rect 1010 440 1062 492
rect 814 346 866 398
rect 900 -382 952 -330
rect 1290 440 1342 492
rect 1094 346 1146 398
rect 1180 -382 1232 -330
rect 1570 440 1622 492
rect 1374 346 1426 398
rect 1460 -382 1512 -330
rect 1850 440 1902 492
rect 1654 346 1706 398
rect 1740 -382 1792 -330
rect 2130 440 2182 492
rect 1934 346 1986 398
rect 2020 -382 2072 -330
rect 2410 440 2462 492
rect 2214 346 2266 398
rect 2300 -382 2352 -330
rect 2690 440 2742 492
rect 2494 346 2546 398
rect 2580 -382 2632 -330
rect 2970 440 3022 492
rect 2774 346 2826 398
rect 2860 -382 2912 -330
rect 3238 238 3290 290
rect 3140 -382 3192 -330
rect 254 -1114 306 -1062
rect 534 -1114 586 -1062
rect 814 -1114 866 -1062
rect 1094 -1114 1146 -1062
rect 1934 -1114 1986 -1062
rect 2214 -1114 2266 -1062
rect 2494 -1114 2546 -1062
rect 2774 -1114 2826 -1062
rect 3054 -1114 3106 -1062
rect 1374 -1230 1426 -1178
rect 1654 -1230 1706 -1178
rect 414 -1514 466 -1462
rect 2478 -1424 2530 -1372
rect 890 -1876 942 -1824
rect 2774 -1876 2826 -1824
rect 330 -1964 382 -1912
rect 610 -1964 662 -1912
rect 178 -2064 230 -2012
rect 254 -2164 306 -2112
rect 458 -2064 510 -2012
rect 534 -2164 586 -2112
rect 814 -2164 866 -2112
rect 1450 -1964 1502 -1912
rect 1730 -1964 1782 -1912
rect 2570 -1964 2622 -1912
rect 1298 -2064 1350 -2012
rect 1094 -2164 1146 -2112
rect 1374 -2164 1426 -2112
rect 1578 -2064 1630 -2012
rect 1654 -2164 1706 -2112
rect 2418 -2064 2470 -2012
rect 1934 -2164 1986 -2112
rect 2214 -2164 2266 -2112
rect 2494 -2164 2546 -2112
rect 2698 -2064 2750 -2012
rect 2850 -1964 2902 -1912
rect 2774 -2164 2826 -2112
rect 178 -2888 230 -2836
rect 458 -2888 510 -2836
rect 738 -2884 790 -2832
rect 330 -2988 382 -2936
rect 1018 -2884 1070 -2832
rect 1298 -2888 1350 -2836
rect 1578 -2888 1630 -2836
rect 1858 -2884 1910 -2832
rect 610 -2988 662 -2936
rect 890 -2988 942 -2936
rect 1170 -2988 1222 -2936
rect 1450 -2988 1502 -2936
rect 254 -3708 306 -3656
rect 534 -3708 586 -3656
rect 814 -3708 866 -3656
rect 890 -3808 942 -3756
rect 1094 -3708 1146 -3656
rect 1374 -3708 1426 -3656
rect 1170 -3808 1222 -3756
rect 738 -3908 790 -3856
rect 1018 -3908 1070 -3856
rect 2138 -2884 2190 -2832
rect 2418 -2888 2470 -2836
rect 2698 -2888 2750 -2836
rect 1730 -2988 1782 -2936
rect 2010 -2988 2062 -2936
rect 2290 -2988 2342 -2936
rect 2570 -2988 2622 -2936
rect 2850 -2988 2902 -2936
rect 1654 -3708 1706 -3656
rect 1934 -3708 1986 -3656
rect 2010 -3808 2062 -3756
rect 1858 -3908 1910 -3856
rect 2214 -3708 2266 -3656
rect 2494 -3708 2546 -3656
rect 2774 -3708 2826 -3656
rect 2290 -3808 2342 -3756
rect 2138 -3908 2190 -3856
rect 1458 -4170 1510 -4118
rect 1578 -4262 1630 -4210
rect 1374 -4986 1426 -4934
rect 1654 -4986 1706 -4934
rect 1296 -5090 1348 -5038
rect 1458 -5170 1510 -5118
rect 1820 -4170 1872 -4118
rect 1734 -5076 1786 -5024
rect 1576 -5780 1628 -5728
rect 1330 -5876 1382 -5824
<< metal2 >>
rect -390 1016 210 1026
rect -390 706 210 716
rect 3028 1016 3628 1026
rect 3028 706 3628 716
rect -120 440 -110 492
rect -58 440 170 492
rect 222 440 450 492
rect 502 440 730 492
rect 782 440 1010 492
rect 1062 440 1290 492
rect 1342 440 1570 492
rect 1622 440 1850 492
rect 1902 440 2130 492
rect 2182 440 2410 492
rect 2462 440 2690 492
rect 2742 440 2970 492
rect 3022 440 3032 492
rect -190 346 -26 398
rect 26 346 36 398
rect 244 346 254 398
rect 306 396 316 398
rect 524 396 534 398
rect 306 346 534 396
rect 586 396 596 398
rect 804 396 814 398
rect 586 346 814 396
rect 866 396 876 398
rect 1084 396 1094 398
rect 866 346 1094 396
rect 1146 396 1156 398
rect 1364 396 1374 398
rect 1146 346 1374 396
rect 1426 396 1436 398
rect 1644 396 1654 398
rect 1426 346 1654 396
rect 1706 396 1716 398
rect 1924 396 1934 398
rect 1706 346 1934 396
rect 1986 396 1996 398
rect 2204 396 2214 398
rect 1986 346 2214 396
rect 2266 396 2276 398
rect 2484 396 2494 398
rect 2266 346 2494 396
rect 2546 396 2556 398
rect 2764 396 2774 398
rect 2546 346 2774 396
rect 2826 396 2836 398
rect 3338 396 3390 398
rect 2826 346 3390 396
rect -190 -1178 -138 346
rect 3238 290 3290 300
rect 50 -382 60 -330
rect 112 -382 340 -330
rect 392 -382 620 -330
rect 672 -382 900 -330
rect 952 -382 1180 -330
rect 1232 -382 1460 -330
rect 1512 -382 1522 -330
rect 1730 -382 1740 -330
rect 1792 -382 2020 -330
rect 2072 -382 2300 -330
rect 2352 -382 2580 -330
rect 2632 -382 2860 -330
rect 2912 -382 3140 -330
rect 3192 -382 3202 -330
rect -36 -1114 -26 -1062
rect 26 -1114 254 -1062
rect 306 -1114 534 -1062
rect 586 -1114 814 -1062
rect 866 -1114 1094 -1062
rect 1146 -1114 1934 -1062
rect 1986 -1114 2214 -1062
rect 2266 -1114 2494 -1062
rect 2546 -1114 2774 -1062
rect 2826 -1114 3054 -1062
rect 3106 -1114 3116 -1062
rect -190 -1230 1374 -1178
rect 1426 -1230 1436 -1178
rect 414 -1462 466 -1452
rect 414 -1824 466 -1514
rect 964 -1466 1016 -1230
rect 1514 -1258 1566 -1114
rect 3238 -1178 3290 238
rect 1644 -1230 1654 -1178
rect 1706 -1230 3290 -1178
rect 3338 -1258 3390 346
rect 1514 -1310 3390 -1258
rect 2478 -1372 2530 -1362
rect 1954 -1466 2000 -1464
rect 2478 -1466 2530 -1424
rect 964 -1518 2530 -1466
rect 414 -1876 890 -1824
rect 942 -1876 952 -1824
rect 1954 -1912 2000 -1518
rect 2916 -1824 2972 -1310
rect 2764 -1876 2774 -1824
rect 2826 -1876 2972 -1824
rect 2916 -1878 2972 -1876
rect 320 -1964 330 -1912
rect 382 -1964 610 -1912
rect 662 -1964 1450 -1912
rect 1502 -1964 1730 -1912
rect 1782 -1964 2570 -1912
rect 2622 -1964 2850 -1912
rect 2902 -1964 3104 -1912
rect -76 -2064 178 -2012
rect 230 -2064 458 -2012
rect 510 -2064 1298 -2012
rect 1350 -2064 1578 -2012
rect 1630 -2064 2418 -2012
rect 2470 -2064 2698 -2012
rect 2750 -2064 2760 -2012
rect -76 -3856 -24 -2064
rect 58 -2164 254 -2112
rect 306 -2164 534 -2112
rect 586 -2164 814 -2112
rect 866 -2164 1094 -2112
rect 1146 -2164 1374 -2112
rect 1426 -2164 1654 -2112
rect 1706 -2164 1934 -2112
rect 1986 -2164 2214 -2112
rect 2266 -2164 2494 -2112
rect 2546 -2164 2774 -2112
rect 2826 -2164 3022 -2112
rect 58 -3656 110 -2164
rect 728 -2836 738 -2832
rect 168 -2888 178 -2836
rect 230 -2888 458 -2836
rect 510 -2884 738 -2836
rect 790 -2836 800 -2832
rect 1008 -2836 1018 -2832
rect 790 -2884 1018 -2836
rect 1070 -2836 1080 -2832
rect 1848 -2836 1858 -2832
rect 1070 -2884 1298 -2836
rect 510 -2888 1298 -2884
rect 1350 -2888 1578 -2836
rect 1630 -2884 1858 -2836
rect 1910 -2836 1920 -2832
rect 2128 -2836 2138 -2832
rect 1910 -2884 2138 -2836
rect 2190 -2836 2200 -2832
rect 2190 -2884 2418 -2836
rect 1630 -2888 2418 -2884
rect 2470 -2888 2698 -2836
rect 2750 -2888 2760 -2836
rect 320 -2988 330 -2936
rect 382 -2988 610 -2936
rect 662 -2988 890 -2936
rect 942 -2988 1170 -2936
rect 1222 -2988 1450 -2936
rect 1502 -2988 1730 -2936
rect 1782 -2988 2010 -2936
rect 2062 -2988 2290 -2936
rect 2342 -2988 2570 -2936
rect 2622 -2988 2850 -2936
rect 2902 -2988 2912 -2936
rect 330 -2990 2902 -2988
rect 2970 -3656 3022 -2164
rect 58 -3708 254 -3656
rect 306 -3708 534 -3656
rect 586 -3708 814 -3656
rect 866 -3708 1094 -3656
rect 1146 -3708 1374 -3656
rect 1426 -3708 1654 -3656
rect 1706 -3708 1934 -3656
rect 1986 -3708 2214 -3656
rect 2266 -3708 2494 -3656
rect 2546 -3708 2774 -3656
rect 2826 -3708 3022 -3656
rect 3052 -3756 3104 -1964
rect 880 -3808 890 -3756
rect 942 -3808 1170 -3756
rect 1222 -3808 2010 -3756
rect 2062 -3808 2290 -3756
rect 2342 -3808 3104 -3756
rect -76 -3908 738 -3856
rect 790 -3908 1018 -3856
rect 1070 -3908 1858 -3856
rect 1910 -3908 2138 -3856
rect 2190 -3908 2200 -3856
rect 1448 -4170 1458 -4118
rect 1510 -4170 1820 -4118
rect 1872 -4170 1882 -4118
rect 1568 -4262 1578 -4210
rect 1630 -4262 1876 -4210
rect 1364 -4986 1374 -4934
rect 1426 -4986 1654 -4934
rect 1706 -4986 1716 -4934
rect 1724 -5036 1734 -5024
rect 1286 -5090 1296 -5038
rect 1348 -5090 1358 -5038
rect 1554 -5070 1734 -5036
rect 1296 -5728 1348 -5090
rect 1554 -5118 1588 -5070
rect 1724 -5076 1734 -5070
rect 1786 -5076 1796 -5024
rect 1448 -5170 1458 -5118
rect 1510 -5170 1588 -5118
rect 1296 -5780 1576 -5728
rect 1628 -5780 1638 -5728
rect 1826 -5824 1876 -4262
rect 1320 -5876 1330 -5824
rect 1382 -5876 1876 -5824
<< via2 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
<< metal3 >>
rect -400 1016 220 1021
rect -400 716 -390 1016
rect 210 716 220 1016
rect -400 711 220 716
rect 3018 1016 3638 1021
rect 3018 716 3028 1016
rect 3628 716 3638 1016
rect 3018 711 3638 716
<< via3 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
<< metal4 >>
rect -391 1016 211 1017
rect -391 716 -390 1016
rect 210 716 211 1016
rect -391 715 211 716
rect 3027 1016 3629 1017
rect 3027 716 3028 1016
rect 3628 716 3629 1016
rect 3027 715 3629 716
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm1
timestamp 1732509526
transform 1 0 0 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm2
timestamp 1732509526
transform 1 0 280 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm3
timestamp 1732509526
transform 1 0 560 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm4
timestamp 1732509526
transform 1 0 840 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm5
timestamp 1732509526
transform 1 0 1120 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm6
timestamp 1732509526
transform 1 0 1400 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm7
timestamp 1732509526
transform 1 0 1680 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm8
timestamp 1732509526
transform 1 0 1960 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm9
timestamp 1732509526
transform 1 0 2240 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm10
timestamp 1732509526
transform 1 0 2520 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm11
timestamp 1732509526
transform 1 0 2800 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm12
timestamp 1732509526
transform 1 0 3080 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm13
timestamp 1732509526
transform 1 0 0 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm14
timestamp 1732509526
transform 1 0 280 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm15
timestamp 1732509526
transform 1 0 560 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm16
timestamp 1732509526
transform 1 0 840 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm17
timestamp 1732509526
transform 1 0 1120 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm18
timestamp 1732509526
transform 1 0 1400 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm19
timestamp 1732509526
transform 1 0 1680 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm20
timestamp 1732509526
transform 1 0 1960 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm21
timestamp 1732509526
transform 1 0 2240 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm22
timestamp 1732509526
transform 1 0 2520 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm23
timestamp 1732509526
transform 1 0 2800 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm24
timestamp 1732509526
transform 1 0 3080 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__nfet_01v8_PHZV97  xm25
timestamp 1732509526
transform 1 0 280 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm26
timestamp 1732509526
transform 1 0 560 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm27
timestamp 1732509526
transform 1 0 840 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm28
timestamp 1732509526
transform 1 0 1120 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm29
timestamp 1732509526
transform 1 0 1400 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm30
timestamp 1732509526
transform 1 0 1680 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm31
timestamp 1732509526
transform 1 0 1960 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm32
timestamp 1732509526
transform 1 0 2240 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm33
timestamp 1732509526
transform 1 0 2520 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm34
timestamp 1732509526
transform 1 0 2800 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm35
timestamp 1732509526
transform 1 0 280 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm36
timestamp 1732509526
transform 1 0 560 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm37
timestamp 1732509526
transform 1 0 840 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm38
timestamp 1732509526
transform 1 0 1120 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm39
timestamp 1732509526
transform 1 0 1400 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm40
timestamp 1732509526
transform 1 0 1680 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm41
timestamp 1732509526
transform 1 0 1960 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm42
timestamp 1732509526
transform 1 0 2240 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm43
timestamp 1732509526
transform 1 0 2520 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm44
timestamp 1732509526
transform 1 0 2800 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm45
timestamp 1732509526
transform 1 0 1400 0 1 -4600
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm46
timestamp 1732509526
transform 1 0 1680 0 1 -4600
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_72KZQ8  xm47
timestamp 1732423020
transform 1 0 1399 0 1 -5427
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm48
timestamp 1732423020
transform 1 0 1679 0 1 -5427
box -73 -257 73 257
<< labels >>
rlabel metal1 -1936 -1298 -1836 -1198 1 M5_net
port 2 n
rlabel metal1 -1946 -1568 -1846 -1468 1 CLK
port 3 n
rlabel metal1 -1942 -1838 -1842 -1738 1 M6_net
port 4 n
rlabel metal1 706 670 806 770 1 VDD
port 1 n
<< properties >>
string FIXED_BBOX -446 -1652 3684 1072
<< end >>
