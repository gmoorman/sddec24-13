magic
tech sky130B
magscale 1 2
timestamp 1731394619
<< nwell >>
rect -374 -1780 3012 1200
<< mvnsubdiff >>
rect -308 1122 2946 1134
rect -308 1022 -134 1122
rect 2772 1022 2946 1122
rect -308 1010 2946 1022
rect -308 960 -184 1010
rect -308 -1540 -296 960
rect -196 -1540 -184 960
rect -308 -1590 -184 -1540
rect 2822 960 2946 1010
rect 2822 -1540 2834 960
rect 2934 -1540 2946 960
rect 2822 -1590 2946 -1540
rect -308 -1602 2946 -1590
rect -308 -1702 -134 -1602
rect 2772 -1702 2946 -1602
rect -308 -1714 2946 -1702
<< mvnsubdiffcont >>
rect -134 1022 2772 1122
rect -296 -1540 -196 960
rect 2834 -1540 2934 960
rect -134 -1702 2772 -1602
<< locali >>
rect -296 960 -196 1122
rect -296 -1702 -196 -1540
rect 2834 960 2934 1122
rect 2834 -1702 2934 -1540
<< viali >>
rect -196 1022 -134 1122
rect -134 1022 2772 1122
rect 2772 1022 2834 1122
rect -296 -1471 -196 891
rect 2834 -1471 2934 891
rect -196 -1702 -134 -1602
rect -134 -1702 2772 -1602
rect 2772 -1702 2834 -1602
<< metal1 >>
rect -302 1122 2940 1128
rect -302 1022 -196 1122
rect 2834 1022 2940 1122
rect -302 1016 2940 1022
rect -302 891 -190 1016
rect -302 -1471 -296 891
rect -196 -1471 -190 891
rect 410 716 420 1016
rect 730 822 782 1016
rect 700 722 800 822
rect -110 492 -58 502
rect -110 -684 -58 440
rect 170 492 222 502
rect -26 398 26 408
rect -26 336 26 346
rect -18 246 18 336
rect -18 -308 18 -246
rect 60 -330 112 -30
rect -18 -470 18 -408
rect -18 -1052 18 -962
rect -26 -1062 26 -1052
rect -26 -1124 26 -1114
rect 60 -1178 112 -382
rect 170 -684 222 440
rect 450 492 502 502
rect 254 398 306 408
rect 254 336 306 346
rect 262 246 298 336
rect 262 -308 298 -246
rect 340 -330 392 -30
rect 262 -470 298 -408
rect 340 -682 392 -382
rect 450 -684 502 440
rect 730 492 782 722
rect 2218 716 2228 1016
rect 2828 891 2940 1016
rect 534 398 586 408
rect 534 336 586 346
rect 542 246 578 336
rect 542 -308 578 -246
rect 620 -330 672 -30
rect 542 -470 578 -408
rect 620 -682 672 -382
rect 730 -684 782 440
rect 1010 492 1062 502
rect 814 398 866 408
rect 814 336 866 346
rect 822 246 858 336
rect 822 -308 858 -246
rect 900 -330 952 -30
rect 822 -470 858 -408
rect 900 -682 952 -382
rect 1010 -684 1062 440
rect 1290 492 1342 502
rect 1094 398 1146 408
rect 1094 336 1146 346
rect 1102 246 1138 336
rect 1102 -308 1138 -246
rect 1180 -330 1232 -30
rect 1102 -470 1138 -408
rect 1180 -682 1232 -382
rect 1290 -684 1342 440
rect 1570 492 1622 502
rect 1374 398 1426 408
rect 1374 336 1426 346
rect 1382 246 1418 336
rect 1382 -308 1418 -246
rect 1460 -330 1512 -30
rect 1382 -470 1418 -408
rect 1460 -682 1512 -382
rect 1570 -684 1622 440
rect 1850 492 1902 502
rect 1654 398 1706 408
rect 1654 336 1706 346
rect 1662 246 1698 336
rect 1662 -308 1698 -246
rect 1740 -330 1792 -30
rect 1662 -470 1698 -408
rect 1740 -682 1792 -382
rect 1850 -684 1902 440
rect 2130 492 2182 502
rect 1934 398 1986 408
rect 1934 336 1986 346
rect 1942 246 1978 336
rect 1942 -308 1978 -246
rect 2020 -330 2072 -30
rect 1942 -470 1978 -408
rect 2020 -682 2072 -382
rect 2130 -684 2182 440
rect 2410 492 2462 502
rect 2214 398 2266 408
rect 2214 336 2266 346
rect 2222 246 2258 336
rect 2222 -308 2258 -246
rect 2300 -330 2352 -30
rect 2222 -470 2258 -408
rect 2300 -682 2352 -382
rect 2410 -684 2462 440
rect 2668 282 2678 290
rect 2502 246 2678 282
rect 2668 238 2678 246
rect 2730 238 2740 290
rect 2502 -308 2538 -246
rect 2580 -330 2632 -30
rect 2502 -470 2538 -408
rect 262 -1052 298 -962
rect 542 -1052 578 -962
rect 822 -1052 858 -962
rect 254 -1062 306 -1052
rect 254 -1124 306 -1114
rect 534 -1062 586 -1052
rect 534 -1124 586 -1114
rect 814 -1062 866 -1052
rect 814 -1124 866 -1114
rect 1102 -1168 1138 -962
rect 1382 -1168 1418 -962
rect 1662 -1052 1698 -962
rect 1942 -1052 1978 -962
rect 2222 -1052 2258 -962
rect 2502 -1052 2538 -962
rect 1654 -1062 1706 -1052
rect 1654 -1124 1706 -1114
rect 1934 -1062 1986 -1052
rect 1934 -1124 1986 -1114
rect 2214 -1062 2266 -1052
rect 2214 -1124 2266 -1114
rect 2494 -1062 2546 -1052
rect 2494 -1124 2546 -1114
rect 2580 -1160 2632 -382
rect 1094 -1178 1146 -1168
rect 50 -1230 60 -1178
rect 112 -1230 122 -1178
rect 60 -1324 112 -1230
rect 1094 -1240 1146 -1230
rect 1374 -1178 1426 -1168
rect 1374 -1240 1426 -1230
rect 1124 -1320 1224 -1284
rect 22 -1424 122 -1324
rect 1124 -1372 1234 -1320
rect 1286 -1372 1296 -1320
rect 1124 -1384 1224 -1372
rect 2580 -1384 2632 -1212
rect -302 -1596 -190 -1471
rect 2564 -1484 2664 -1384
rect 2828 -1471 2834 891
rect 2934 -1471 2940 891
rect 2828 -1596 2940 -1471
rect -302 -1602 2940 -1596
rect -302 -1702 -196 -1602
rect 2834 -1702 2940 -1602
rect -302 -1708 2940 -1702
<< via1 >>
rect -190 716 410 1016
rect -110 440 -58 492
rect 170 440 222 492
rect -26 346 26 398
rect 60 -382 112 -330
rect -26 -1114 26 -1062
rect 450 440 502 492
rect 254 346 306 398
rect 340 -382 392 -330
rect 2228 716 2828 1016
rect 730 440 782 492
rect 534 346 586 398
rect 620 -382 672 -330
rect 1010 440 1062 492
rect 814 346 866 398
rect 900 -382 952 -330
rect 1290 440 1342 492
rect 1094 346 1146 398
rect 1180 -382 1232 -330
rect 1570 440 1622 492
rect 1374 346 1426 398
rect 1460 -382 1512 -330
rect 1850 440 1902 492
rect 1654 346 1706 398
rect 1740 -382 1792 -330
rect 2130 440 2182 492
rect 1934 346 1986 398
rect 2020 -382 2072 -330
rect 2410 440 2462 492
rect 2214 346 2266 398
rect 2300 -382 2352 -330
rect 2678 238 2730 290
rect 2580 -382 2632 -330
rect 254 -1114 306 -1062
rect 534 -1114 586 -1062
rect 814 -1114 866 -1062
rect 1654 -1114 1706 -1062
rect 1934 -1114 1986 -1062
rect 2214 -1114 2266 -1062
rect 2494 -1114 2546 -1062
rect 60 -1230 112 -1178
rect 1094 -1230 1146 -1178
rect 1374 -1230 1426 -1178
rect 2580 -1212 2632 -1160
rect 1234 -1372 1286 -1320
<< metal2 >>
rect -190 1016 410 1026
rect -190 706 410 716
rect 2228 1016 2828 1026
rect 2228 706 2828 716
rect -120 440 -110 492
rect -58 440 170 492
rect 222 440 450 492
rect 502 440 730 492
rect 782 440 1010 492
rect 1062 440 1290 492
rect 1342 440 1570 492
rect 1622 440 1850 492
rect 1902 440 2130 492
rect 2182 440 2410 492
rect 2462 440 2472 492
rect -190 346 -26 398
rect 26 346 36 398
rect 244 346 254 398
rect 306 346 534 398
rect 586 346 814 398
rect 866 346 1094 398
rect 1146 346 1374 398
rect 1426 346 1654 398
rect 1706 346 1934 398
rect 1986 346 2214 398
rect 2266 346 2826 398
rect -190 -1178 -138 346
rect 244 344 2826 346
rect 2678 290 2730 300
rect 50 -382 60 -330
rect 112 -382 340 -330
rect 392 -382 620 -330
rect 672 -382 900 -330
rect 952 -382 1180 -330
rect 1232 -382 1242 -330
rect 1450 -382 1460 -330
rect 1512 -382 1740 -330
rect 1792 -382 2020 -330
rect 2072 -382 2300 -330
rect 2352 -382 2580 -330
rect 2632 -382 2642 -330
rect -36 -1114 -26 -1062
rect 26 -1114 254 -1062
rect 306 -1114 534 -1062
rect 586 -1114 814 -1062
rect 866 -1114 1654 -1062
rect 1706 -1114 1934 -1062
rect 1986 -1114 2214 -1062
rect 2266 -1114 2494 -1062
rect 2546 -1114 2556 -1062
rect 60 -1178 112 -1168
rect -190 -1230 60 -1178
rect 112 -1230 1094 -1178
rect 1146 -1230 1156 -1178
rect 60 -1240 112 -1230
rect 1234 -1258 1286 -1114
rect 2570 -1178 2580 -1160
rect 1364 -1230 1374 -1178
rect 1426 -1212 2580 -1178
rect 2632 -1178 2642 -1160
rect 2678 -1178 2730 238
rect 2632 -1212 2730 -1178
rect 1426 -1230 2730 -1212
rect 2774 -1258 2826 344
rect 1234 -1310 2826 -1258
rect 1234 -1320 1286 -1310
rect 1234 -1382 1286 -1372
<< via2 >>
rect -190 716 410 1016
rect 2228 716 2828 1016
<< metal3 >>
rect -200 1016 420 1021
rect -200 716 -190 1016
rect 410 716 420 1016
rect -200 711 420 716
rect 2218 1016 2838 1021
rect 2218 716 2228 1016
rect 2828 716 2838 1016
rect 2218 711 2838 716
<< via3 >>
rect -190 716 410 1016
rect 2228 716 2828 1016
<< metal4 >>
rect -191 1016 411 1017
rect -191 716 -190 1016
rect 410 716 411 1016
rect -191 715 411 716
rect 2227 1016 2829 1017
rect 2227 716 2228 1016
rect 2828 716 2829 1016
rect 2227 715 2829 716
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm1
timestamp 1731387447
transform 1 0 0 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm2
timestamp 1731387447
transform 1 0 280 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm3
timestamp 1731387447
transform 1 0 560 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm4
timestamp 1731387447
transform 1 0 840 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm5
timestamp 1731387447
transform 1 0 1120 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm6
timestamp 1731387447
transform 1 0 1400 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm7
timestamp 1731387447
transform 1 0 1680 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm8
timestamp 1731387447
transform 1 0 1960 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm9
timestamp 1731387447
transform 1 0 2240 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm10
timestamp 1731387447
transform 1 0 2520 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm11
timestamp 1731387447
transform 1 0 0 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm12
timestamp 1731387447
transform 1 0 280 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm13
timestamp 1731387447
transform 1 0 560 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm14
timestamp 1731387447
transform 1 0 840 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm15
timestamp 1731387447
transform 1 0 1120 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm16
timestamp 1731387447
transform 1 0 1400 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm17
timestamp 1731387447
transform 1 0 1680 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm18
timestamp 1731387447
transform 1 0 1960 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm19
timestamp 1731387447
transform 1 0 2240 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm20
timestamp 1731387447
transform 1 0 2520 0 1 -716
box -109 -300 109 300
<< labels >>
rlabel metal1 2564 -1484 2664 -1384 1 M6_net
port 3 n
rlabel metal1 1124 -1384 1224 -1284 1 CLK
port 1 n
rlabel metal1 700 722 800 822 1 VDD
port 4 n
rlabel metal1 22 -1424 122 -1324 1 M5_net
port 2 n
<< properties >>
string FIXED_BBOX -246 -1652 2884 1072
<< end >>
