* NGSPICE file created from 4x4crossbar.ext - technology: sky130B

.subckt sky130_fd_pr_reram__reram_cell_X TE BE
X0 TE BE sky130_fd_pr_reram__reram_cell area_ox=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B a_50_n700# a_n242_n922# a_n108_n700# a_n50_n788#
X0 a_50_n700# a_n50_n788# a_n108_n700# a_n242_n922# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=0.5
.ends

.subckt x1T1R SL VSS WL BL
XXR1 BL XR1/BE sky130_fd_pr_reram__reram_cell_X
XXM1 XR1/BE VSS SL WL sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
.ends

.subckt x2x2crossbar BL2 WL2 WL1 BL1 VSS SL2 SL1
Xx1 SL1 VSS WL1 BL1 x1T1R
Xx2 SL2 VSS WL1 BL2 x1T1R
Xx3 SL1 VSS WL2 BL1 x1T1R
Xx4 SL2 VSS WL2 BL2 x1T1R
.ends

.subckt x4x4crossbar BL1 BL2 SL2 SL1 BL3 BL4 SL4 SL3 WL2 WL1 WL4 WL3 VSS
Xx1 BL2 WL2 WL1 BL1 VSS SL2 SL1 x2x2crossbar
Xx3 BL4 WL2 WL1 BL3 VSS SL4 SL3 x2x2crossbar
Xx2 BL2 WL4 WL3 BL1 VSS SL2 SL1 x2x2crossbar
Xx4 BL4 WL4 WL3 BL3 VSS SL4 SL3 x2x2crossbar
.ends

