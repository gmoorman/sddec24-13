magic
tech sky130B
magscale 1 2
timestamp 1733700048
<< nwell >>
rect -296 -2137 296 2137
<< pmoslvt >>
rect -100 118 100 1918
rect -100 -1918 100 -118
<< pdiff >>
rect -158 1906 -100 1918
rect -158 130 -146 1906
rect -112 130 -100 1906
rect -158 118 -100 130
rect 100 1906 158 1918
rect 100 130 112 1906
rect 146 130 158 1906
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -1906 -146 -130
rect -112 -1906 -100 -130
rect -158 -1918 -100 -1906
rect 100 -130 158 -118
rect 100 -1906 112 -130
rect 146 -1906 158 -130
rect 100 -1918 158 -1906
<< pdiffc >>
rect -146 130 -112 1906
rect 112 130 146 1906
rect -146 -1906 -112 -130
rect 112 -1906 146 -130
<< nsubdiff >>
rect -260 2067 -164 2101
rect 164 2067 260 2101
rect -260 2005 -226 2067
rect 226 2005 260 2067
rect -260 -2067 -226 -2005
rect 226 -2067 260 -2005
rect -260 -2101 -164 -2067
rect 164 -2101 260 -2067
<< nsubdiffcont >>
rect -164 2067 164 2101
rect -260 -2005 -226 2005
rect 226 -2005 260 2005
rect -164 -2101 164 -2067
<< poly >>
rect -100 1999 100 2015
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -100 1918 100 1965
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -1965 100 -1918
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -100 -2015 100 -1999
<< polycont >>
rect -84 1965 84 1999
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1999 84 -1965
<< locali >>
rect -260 2067 -164 2101
rect 164 2067 260 2101
rect -260 2005 -226 2067
rect 226 2005 260 2067
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -146 1906 -112 1922
rect -146 114 -112 130
rect 112 1906 146 1922
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -1922 -112 -1906
rect 112 -130 146 -114
rect 112 -1922 146 -1906
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -260 -2067 -226 -2005
rect 226 -2067 260 -2005
rect -260 -2101 -164 -2067
rect 164 -2101 260 -2067
<< viali >>
rect -84 1965 84 1999
rect -146 130 -112 1906
rect 112 130 146 1906
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1906 -112 -130
rect 112 -1906 146 -130
rect -84 -1999 84 -1965
<< metal1 >>
rect -96 1999 96 2005
rect -96 1965 -84 1999
rect 84 1965 96 1999
rect -96 1959 96 1965
rect -152 1906 -106 1918
rect -152 130 -146 1906
rect -112 130 -106 1906
rect -152 118 -106 130
rect 106 1906 152 1918
rect 106 130 112 1906
rect 146 130 152 1906
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -1906 -146 -130
rect -112 -1906 -106 -130
rect -152 -1918 -106 -1906
rect 106 -130 152 -118
rect 106 -1906 112 -130
rect 146 -1906 152 -130
rect 106 -1918 152 -1906
rect -96 -1965 96 -1959
rect -96 -1999 -84 -1965
rect 84 -1999 96 -1965
rect -96 -2005 96 -1999
<< properties >>
string FIXED_BBOX -243 -2084 243 2084
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 9.0 l 1.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
