magic
tech sky130B
magscale 1 2
timestamp 1733216309
<< error_p >>
rect -29 241 29 247
rect -29 207 -17 241
rect -29 201 29 207
<< pwell >>
rect -99 -257 99 195
<< nmos >>
rect -15 -231 15 169
<< ndiff >>
rect -73 156 -15 169
rect -73 122 -61 156
rect -27 122 -15 156
rect -73 88 -15 122
rect -73 54 -61 88
rect -27 54 -15 88
rect -73 20 -15 54
rect -73 -14 -61 20
rect -27 -14 -15 20
rect -73 -48 -15 -14
rect -73 -82 -61 -48
rect -27 -82 -15 -48
rect -73 -116 -15 -82
rect -73 -150 -61 -116
rect -27 -150 -15 -116
rect -73 -184 -15 -150
rect -73 -218 -61 -184
rect -27 -218 -15 -184
rect -73 -231 -15 -218
rect 15 156 73 169
rect 15 122 27 156
rect 61 122 73 156
rect 15 88 73 122
rect 15 54 27 88
rect 61 54 73 88
rect 15 20 73 54
rect 15 -14 27 20
rect 61 -14 73 20
rect 15 -48 73 -14
rect 15 -82 27 -48
rect 61 -82 73 -48
rect 15 -116 73 -82
rect 15 -150 27 -116
rect 61 -150 73 -116
rect 15 -184 73 -150
rect 15 -218 27 -184
rect 61 -218 73 -184
rect 15 -231 73 -218
<< ndiffc >>
rect -61 122 -27 156
rect -61 54 -27 88
rect -61 -14 -27 20
rect -61 -82 -27 -48
rect -61 -150 -27 -116
rect -61 -218 -27 -184
rect 27 122 61 156
rect 27 54 61 88
rect 27 -14 61 20
rect 27 -82 61 -48
rect 27 -150 61 -116
rect 27 -218 61 -184
<< poly >>
rect -33 241 33 257
rect -33 207 -17 241
rect 17 207 33 241
rect -33 191 33 207
rect -15 169 15 191
rect -15 -257 15 -231
<< polycont >>
rect -17 207 17 241
<< locali >>
rect -33 207 -17 241
rect 17 207 33 241
rect -61 156 -27 173
rect -61 88 -27 96
rect -61 20 -27 24
rect -61 -86 -27 -82
rect -61 -158 -27 -150
rect -61 -235 -27 -218
rect 27 156 61 173
rect 27 88 61 96
rect 27 20 61 24
rect 27 -86 61 -82
rect 27 -158 61 -150
rect 27 -235 61 -218
<< viali >>
rect -17 207 17 241
rect -61 122 -27 130
rect -61 96 -27 122
rect -61 54 -27 58
rect -61 24 -27 54
rect -61 -48 -27 -14
rect -61 -116 -27 -86
rect -61 -120 -27 -116
rect -61 -184 -27 -158
rect -61 -192 -27 -184
rect 27 122 61 130
rect 27 96 61 122
rect 27 54 61 58
rect 27 24 61 54
rect 27 -48 61 -14
rect 27 -116 61 -86
rect 27 -120 61 -116
rect 27 -184 61 -158
rect 27 -192 61 -184
<< metal1 >>
rect -29 241 29 247
rect -29 207 -17 241
rect 17 207 29 241
rect -29 201 29 207
rect -67 130 -21 169
rect -67 96 -61 130
rect -27 96 -21 130
rect -67 58 -21 96
rect -67 24 -61 58
rect -27 24 -21 58
rect -67 -14 -21 24
rect -67 -48 -61 -14
rect -27 -48 -21 -14
rect -67 -86 -21 -48
rect -67 -120 -61 -86
rect -27 -120 -21 -86
rect -67 -158 -21 -120
rect -67 -192 -61 -158
rect -27 -192 -21 -158
rect -67 -231 -21 -192
rect 21 130 67 169
rect 21 96 27 130
rect 61 96 67 130
rect 21 58 67 96
rect 21 24 27 58
rect 61 24 67 58
rect 21 -14 67 24
rect 21 -48 27 -14
rect 61 -48 67 -14
rect 21 -86 67 -48
rect 21 -120 27 -86
rect 61 -120 67 -86
rect 21 -158 67 -120
rect 21 -192 27 -158
rect 61 -192 67 -158
rect 21 -231 67 -192
<< end >>
