magic
tech sky130B
timestamp 1731452249
<< metal1 >>
rect 830 100 1470 200
rect 1150 -1080 1250 100
rect 830 -1180 1470 -1080
<< metal2 >>
rect 680 1170 1460 1270
rect 680 240 1320 340
rect 680 -110 1460 -10
rect 680 -1040 1320 -940
<< metal3 >>
rect 1150 -650 1250 1270
rect 1690 -650 1790 1270
use 1T1R  x1 ~/reram/caravel_user_project_analog/mag
timestamp 1731452249
transform 1 0 860 0 1 -140
box -180 210 395 1415
use 1T1R  x2
timestamp 1731452249
transform 1 0 1400 0 1 -140
box -180 210 395 1415
use 1T1R  x3
timestamp 1731452249
transform 1 0 860 0 1 -1420
box -180 210 395 1415
use 1T1R  x4
timestamp 1731452249
transform 1 0 1400 0 1 -1420
box -180 210 395 1415
<< labels >>
flabel metal2 680 240 780 340 0 FreeSans 128 0 0 0 WL1
port 3 nsew
flabel metal2 680 -1040 780 -940 0 FreeSans 128 0 0 0 WL2
port 4 nsew
flabel metal3 1150 1170 1250 1270 0 FreeSans 128 0 0 0 BL1
port 1 nsew
flabel metal3 1690 1170 1790 1270 0 FreeSans 128 0 0 0 BL2
port 0 nsew
flabel metal1 830 100 930 200 0 FreeSans 128 0 0 0 VSS
port 2 nsew
flabel metal2 680 1170 780 1270 0 FreeSans 128 0 0 0 SL1
port 5 nsew
flabel metal2 680 -110 780 -10 0 FreeSans 128 0 0 0 SL2
port 6 nsew
<< end >>
