** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/8x8.sch
.subckt 8x8 BL1 BL2 BL3 BL4 BL5 BL6 BL7 BL8 SL1 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 SL2 SL3 SL4 SL5 SL6
+ SL7 SL8 VSS
*.PININFO BL1:B BL2:B BL3:B BL4:B BL5:B BL6:B BL7:B BL8:B SL1:B WL1:B WL2:B WL3:B WL4:B WL5:B WL6:B
*+ WL7:B WL8:B SL2:B SL3:B SL4:B SL5:B SL6:B SL7:B SL8:B VSS:B
x1 VSS BL1 BL3 BL2 BL4 SL1 SL2 WL2 WL1 WL4 WL3 SL3 SL4 4x4
x2 VSS BL5 BL7 BL6 BL8 SL1 SL2 WL2 WL1 WL4 WL3 SL3 SL4 4x4
x3 VSS BL5 BL7 BL6 BL8 SL5 SL6 WL6 WL5 WL8 WL7 SL7 SL8 4x4
x4 VSS BL1 BL3 BL2 BL4 SL5 SL6 WL6 WL5 WL8 WL7 SL7 SL8 4x4
.ends

* expanding   symbol:  4x4.sym # of pins=13
** sym_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/4x4.sym
** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/4x4.sch
.subckt 4x4 VSS BL1 BL3 BL2 BL4 SL1 SL2 WL2 WL1 WL4 WL3 SL3 SL4
*.PININFO BL1:B BL2:B SL2:B SL1:B BL3:B BL4:B SL4:B SL3:B WL2:B WL1:B WL4:B WL3:B VSS:B
x1 VSS BL2 BL1 WL1 SL1 WL2 SL2 2x2
x2 VSS BL2 BL1 WL3 SL3 WL4 SL4 2x2
x3 VSS BL4 BL3 WL1 SL1 WL2 SL2 2x2
x4 VSS BL4 BL3 WL3 SL3 WL4 SL4 2x2
.ends


* expanding   symbol:  2x2.sym # of pins=7
** sym_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/2x2.sym
** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/2x2.sch
.subckt 2x2 VSS BL2 BL1 WL1 SL1 WL2 SL2
*.PININFO BL2:B BL1:B VSS:B WL1:B WL2:B SL1:B SL2:B
x1 BL1 WL1 VSS SL1 1T1R
x2 BL2 WL1 VSS SL1 1T1R
x3 BL1 WL2 VSS SL2 1T1R
x4 BL2 WL2 VSS SL2 1T1R
.ends


* expanding   symbol:  1T1R.sym # of pins=4
** sym_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/1T1R.sym
** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/1T1R.sch
.subckt 1T1R BL WL VSS SL
*.PININFO SL:B VSS:B WL:B BL:B
XR1 BL net1 sky130_fd_pr_reram__reram_cell Tfilament_0=3.8e-9 area_ox=1
XM1 net1 WL SL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=1
.ends


.end
