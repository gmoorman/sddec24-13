magic
tech sky130B
timestamp 1733700048
<< pwell >>
rect -148 -814 148 814
<< nmos >>
rect -50 309 50 709
rect -50 -200 50 200
rect -50 -709 50 -309
<< ndiff >>
rect -79 703 -50 709
rect -79 315 -73 703
rect -56 315 -50 703
rect -79 309 -50 315
rect 50 703 79 709
rect 50 315 56 703
rect 73 315 79 703
rect 50 309 79 315
rect -79 194 -50 200
rect -79 -194 -73 194
rect -56 -194 -50 194
rect -79 -200 -50 -194
rect 50 194 79 200
rect 50 -194 56 194
rect 73 -194 79 194
rect 50 -200 79 -194
rect -79 -315 -50 -309
rect -79 -703 -73 -315
rect -56 -703 -50 -315
rect -79 -709 -50 -703
rect 50 -315 79 -309
rect 50 -703 56 -315
rect 73 -703 79 -315
rect 50 -709 79 -703
<< ndiffc >>
rect -73 315 -56 703
rect 56 315 73 703
rect -73 -194 -56 194
rect 56 -194 73 194
rect -73 -703 -56 -315
rect 56 -703 73 -315
<< psubdiff >>
rect -130 779 -82 796
rect 82 779 130 796
rect -130 748 -113 779
rect 113 748 130 779
rect -130 -779 -113 -748
rect 113 -779 130 -748
rect -130 -796 -82 -779
rect 82 -796 130 -779
<< psubdiffcont >>
rect -82 779 82 796
rect -130 -748 -113 748
rect 113 -748 130 748
rect -82 -796 82 -779
<< poly >>
rect -50 745 50 753
rect -50 728 -42 745
rect 42 728 50 745
rect -50 709 50 728
rect -50 290 50 309
rect -50 273 -42 290
rect 42 273 50 290
rect -50 265 50 273
rect -50 236 50 244
rect -50 219 -42 236
rect 42 219 50 236
rect -50 200 50 219
rect -50 -219 50 -200
rect -50 -236 -42 -219
rect 42 -236 50 -219
rect -50 -244 50 -236
rect -50 -273 50 -265
rect -50 -290 -42 -273
rect 42 -290 50 -273
rect -50 -309 50 -290
rect -50 -728 50 -709
rect -50 -745 -42 -728
rect 42 -745 50 -728
rect -50 -753 50 -745
<< polycont >>
rect -42 728 42 745
rect -42 273 42 290
rect -42 219 42 236
rect -42 -236 42 -219
rect -42 -290 42 -273
rect -42 -745 42 -728
<< locali >>
rect -130 779 -82 796
rect 82 779 130 796
rect -130 748 -113 779
rect 113 748 130 779
rect -50 728 -42 745
rect 42 728 50 745
rect -73 703 -56 711
rect -73 307 -56 315
rect 56 703 73 711
rect 56 307 73 315
rect -50 273 -42 290
rect 42 273 50 290
rect -50 219 -42 236
rect 42 219 50 236
rect -73 194 -56 202
rect -73 -202 -56 -194
rect 56 194 73 202
rect 56 -202 73 -194
rect -50 -236 -42 -219
rect 42 -236 50 -219
rect -50 -290 -42 -273
rect 42 -290 50 -273
rect -73 -315 -56 -307
rect -73 -711 -56 -703
rect 56 -315 73 -307
rect 56 -711 73 -703
rect -50 -745 -42 -728
rect 42 -745 50 -728
rect -130 -779 -113 -748
rect 113 -779 130 -748
rect -130 -796 -82 -779
rect 82 -796 130 -779
<< viali >>
rect -42 728 42 745
rect -73 315 -56 703
rect 56 315 73 703
rect -42 273 42 290
rect -42 219 42 236
rect -73 -194 -56 194
rect 56 -194 73 194
rect -42 -236 42 -219
rect -42 -290 42 -273
rect -73 -703 -56 -315
rect 56 -703 73 -315
rect -42 -745 42 -728
<< metal1 >>
rect -48 745 48 748
rect -48 728 -42 745
rect 42 728 48 745
rect -48 725 48 728
rect -76 703 -53 709
rect -76 315 -73 703
rect -56 315 -53 703
rect -76 309 -53 315
rect 53 703 76 709
rect 53 315 56 703
rect 73 315 76 703
rect 53 309 76 315
rect -48 290 48 293
rect -48 273 -42 290
rect 42 273 48 290
rect -48 270 48 273
rect -48 236 48 239
rect -48 219 -42 236
rect 42 219 48 236
rect -48 216 48 219
rect -76 194 -53 200
rect -76 -194 -73 194
rect -56 -194 -53 194
rect -76 -200 -53 -194
rect 53 194 76 200
rect 53 -194 56 194
rect 73 -194 76 194
rect 53 -200 76 -194
rect -48 -219 48 -216
rect -48 -236 -42 -219
rect 42 -236 48 -219
rect -48 -239 48 -236
rect -48 -273 48 -270
rect -48 -290 -42 -273
rect 42 -290 48 -273
rect -48 -293 48 -290
rect -76 -315 -53 -309
rect -76 -703 -73 -315
rect -56 -703 -53 -315
rect -76 -709 -53 -703
rect 53 -315 76 -309
rect 53 -703 56 -315
rect 73 -703 76 -315
rect 53 -709 76 -703
rect -48 -728 48 -725
rect -48 -745 -42 -728
rect 42 -745 48 -728
rect -48 -748 48 -745
<< properties >>
string FIXED_BBOX -121 -787 121 787
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.0 l 1.0 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
