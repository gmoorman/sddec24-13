** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/2x2.sch
.subckt 2x2 BL2 BL1 VSS WL1 WL2 SL1 SL2
*.PININFO BL2:B BL1:B VSS:B WL1:B WL2:B SL1:B SL2:B
x1 BL1 WL1 VSS SL1 1T1R
x2 BL2 WL1 VSS SL1 1T1R
x3 BL1 WL2 VSS SL2 1T1R
x4 BL2 WL2 VSS SL2 1T1R
.ends

* expanding   symbol:  1T1R.sym # of pins=4
** sym_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/1T1R.sym
** sch_path: /home/kivimagi/reram/caravel_user_project_analog/xschem/1T1R.sch
.subckt 1T1R BL WL VSS SL
*.PININFO SL:B VSS:B WL:B BL:B
XR1 BL net1 sky130_fd_pr_reram__reram_cell Tfilament_0=3.8e-9 area_ox=1
XM1 net1 WL SL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 nf=1 m=1
.ends

.end
