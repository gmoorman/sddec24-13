magic
tech sky130B
magscale 1 2
timestamp 1733704917
<< nwell >>
rect -240 -1530 4080 1840
<< pwell >>
rect 4128 -436 4730 1566
<< psubdiff >>
rect 4188 1500 4248 1534
rect 4628 1500 4688 1534
rect 4188 1474 4222 1500
rect 4188 -350 4222 -324
rect 4654 1474 4688 1500
rect 4654 -350 4688 -324
rect 4188 -384 4248 -350
rect 4628 -384 4688 -350
<< mvnsubdiff >>
rect -174 1762 4014 1774
rect -174 1662 0 1762
rect 3840 1662 4014 1762
rect -174 1650 4014 1662
rect -174 1600 -50 1650
rect -174 -1290 -162 1600
rect -62 -1290 -50 1600
rect -174 -1340 -50 -1290
rect 3890 1600 4014 1650
rect 3890 -1290 3902 1600
rect 4002 -1290 4014 1600
rect 3890 -1340 4014 -1290
rect -174 -1352 4014 -1340
rect -174 -1452 0 -1352
rect 3840 -1452 4014 -1352
rect -174 -1464 4014 -1452
<< psubdiffcont >>
rect 4248 1500 4628 1534
rect 4188 -324 4222 1474
rect 4654 -324 4688 1474
rect 4248 -384 4628 -350
<< mvnsubdiffcont >>
rect 0 1662 3840 1762
rect -162 -1290 -62 1600
rect 3902 -1290 4002 1600
rect 0 -1452 3840 -1352
<< locali >>
rect -162 1600 -62 1762
rect -162 -1452 -62 -1290
rect 3902 1600 4002 1762
rect 4188 1500 4248 1534
rect 4628 1500 4688 1534
rect 4188 1474 4222 1500
rect 4188 -350 4222 -324
rect 4654 1474 4688 1500
rect 4654 -350 4688 -324
rect 4188 -384 4248 -350
rect 4628 -384 4688 -350
rect 3902 -1452 4002 -1290
<< viali >>
rect -62 1662 0 1762
rect 0 1662 3840 1762
rect 3840 1662 3902 1762
rect -162 -1201 -62 1511
rect 4406 1534 4468 1538
rect 3902 -1201 4002 1511
rect 4406 1500 4468 1534
rect 4406 1498 4468 1500
rect -62 -1452 0 -1352
rect 0 -1452 3840 -1352
rect 3840 -1452 3902 -1352
<< metal1 >>
rect -168 1762 4008 1768
rect -168 1662 -62 1762
rect 3902 1662 4008 1762
rect -168 1656 4008 1662
rect -168 1511 -56 1656
rect -168 -1201 -162 1511
rect -62 -1201 -56 1511
rect 544 1356 554 1656
rect 3286 1356 3296 1656
rect 3896 1511 4008 1656
rect 1826 1326 1878 1336
rect 1826 1264 1878 1274
rect 1838 1162 1866 1264
rect 98 1126 3610 1162
rect 3652 1068 3680 1356
rect 36 -62 70 92
rect 294 38 328 80
rect 284 28 336 38
rect 284 -34 336 -24
rect 406 -62 440 102
rect 664 38 698 80
rect 654 28 706 38
rect 654 -34 706 -24
rect 778 -62 812 92
rect 1036 38 1070 80
rect 1026 28 1078 38
rect 1026 -34 1078 -24
rect 1148 -62 1182 102
rect 1406 38 1440 80
rect 1396 28 1448 38
rect 1396 -34 1448 -24
rect 1520 -62 1554 92
rect 1778 38 1812 80
rect 1768 28 1820 38
rect 1768 -34 1820 -24
rect 1890 -62 1924 102
rect 2148 38 2182 80
rect 2138 28 2190 38
rect 2138 -34 2190 -24
rect 2262 -62 2296 92
rect 2520 38 2554 80
rect 2510 28 2562 38
rect 2510 -34 2562 -24
rect 2632 -62 2666 102
rect 2890 38 2924 80
rect 2880 28 2932 38
rect 2880 -34 2932 -24
rect 3010 -62 3044 92
rect 3268 38 3302 80
rect 3258 28 3310 38
rect 3258 -34 3310 -24
rect 3380 -62 3414 102
rect 3638 38 3672 80
rect 3628 28 3680 38
rect 3628 -34 3680 -24
rect 36 -92 3820 -62
rect 804 -138 856 -128
rect 804 -200 856 -190
rect 1070 -242 1104 -92
rect 1192 -138 1244 -128
rect 1192 -200 1244 -190
rect 1458 -242 1492 -92
rect 1578 -138 1630 -128
rect 1578 -200 1630 -190
rect 1846 -242 1880 -92
rect 1966 -138 2018 -128
rect 1966 -200 2018 -190
rect 2234 -242 2268 -92
rect 2356 -138 2408 -128
rect 2356 -200 2408 -190
rect 2622 -242 2656 -92
rect 2744 -138 2796 -128
rect 2744 -200 2796 -190
rect 3010 -242 3044 -92
rect 3130 -138 3182 -128
rect 3130 -200 3182 -190
rect 3398 -242 3432 -92
rect 3518 -138 3570 -128
rect 3518 -200 3570 -190
rect 3786 -228 3820 -92
rect -168 -1346 -56 -1201
rect 3896 -1201 3902 1511
rect 4002 -1201 4008 1511
rect 4394 1538 4480 1544
rect 4394 1498 4406 1538
rect 4468 1498 4480 1538
rect 4394 1492 4480 1498
rect 4414 1348 4458 1492
rect 4406 1288 4466 1348
rect 4414 896 4458 1288
rect 4336 866 4540 896
rect 4326 -48 4378 -38
rect 4484 -100 4494 -48
rect 4546 -100 4556 -48
rect 4326 -110 4378 -100
rect 1502 -1246 1512 -1230
rect 872 -1282 1512 -1246
rect 1564 -1246 1574 -1230
rect 3056 -1246 3066 -1230
rect 1564 -1282 2206 -1246
rect 2426 -1282 3066 -1246
rect 3118 -1246 3128 -1230
rect 3118 -1282 3760 -1246
rect 3896 -1346 4008 -1201
rect -168 -1352 4008 -1346
rect -168 -1452 -62 -1352
rect 3902 -1452 4008 -1352
rect -168 -1458 4008 -1452
<< via1 >>
rect -56 1356 544 1656
rect 3296 1356 3896 1656
rect 1826 1274 1878 1326
rect 284 -24 336 28
rect 654 -24 706 28
rect 1026 -24 1078 28
rect 1396 -24 1448 28
rect 1768 -24 1820 28
rect 2138 -24 2190 28
rect 2510 -24 2562 28
rect 2880 -24 2932 28
rect 3258 -24 3310 28
rect 3628 -24 3680 28
rect 804 -190 856 -138
rect 1192 -190 1244 -138
rect 1578 -190 1630 -138
rect 1966 -190 2018 -138
rect 2356 -190 2408 -138
rect 2744 -190 2796 -138
rect 3130 -190 3182 -138
rect 3518 -190 3570 -138
rect 4326 -100 4378 -48
rect 4494 -100 4546 -48
rect 1512 -1282 1564 -1230
rect 3066 -1282 3118 -1230
<< metal2 >>
rect -56 1656 544 1666
rect -56 1346 544 1356
rect 3296 1656 3896 1666
rect 3296 1346 3896 1356
rect 1888 1326 1948 1332
rect 1816 1274 1826 1326
rect 1878 1274 1948 1326
rect 1888 1272 1948 1274
rect 274 -24 284 28
rect 336 -24 654 28
rect 706 -24 1026 28
rect 1078 -24 1396 28
rect 1448 -24 1768 28
rect 1820 -24 2138 28
rect 2190 -24 2510 28
rect 2562 -24 2880 28
rect 2932 -24 3258 28
rect 3310 -24 3628 28
rect 3680 -24 3690 28
rect 4074 -60 4134 -40
rect 4494 -48 4546 -38
rect 4316 -60 4326 -48
rect 2234 -88 4326 -60
rect 794 -190 804 -138
rect 856 -190 1192 -138
rect 1244 -190 1578 -138
rect 1630 -190 1966 -138
rect 2018 -154 2028 -138
rect 2234 -154 2266 -88
rect 4074 -100 4134 -88
rect 4316 -100 4326 -88
rect 4378 -100 4388 -48
rect 2018 -190 2266 -154
rect 2346 -190 2356 -138
rect 2408 -190 2744 -138
rect 2796 -190 3130 -138
rect 3182 -190 3518 -138
rect 3570 -160 3576 -138
rect 4074 -160 4134 -144
rect 4494 -160 4546 -100
rect 3570 -190 4546 -160
rect 4074 -204 4134 -190
rect 1512 -1230 1564 -1220
rect 3066 -1230 3118 -1220
rect 1508 -1342 1568 -1282
rect 3062 -1342 3122 -1282
<< via2 >>
rect -56 1356 544 1656
rect 3296 1356 3896 1656
<< metal3 >>
rect -66 1656 554 1661
rect -66 1356 -56 1656
rect 544 1356 554 1656
rect -66 1351 554 1356
rect 3286 1656 3906 1661
rect 3286 1356 3296 1656
rect 3896 1356 3906 1656
rect 3286 1351 3906 1356
<< via3 >>
rect -56 1356 544 1656
rect 3296 1356 3896 1656
<< metal4 >>
rect -57 1656 545 1657
rect -57 1356 -56 1656
rect 544 1356 545 1656
rect -57 1355 545 1356
rect 3295 1656 3897 1657
rect 3295 1356 3296 1656
rect 3896 1356 3897 1656
rect 3295 1355 3897 1356
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_0
timestamp 1733704561
transform 1 0 958 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_1
timestamp 1733704561
transform 1 0 1346 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_2
timestamp 1733704561
transform 1 0 1734 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_3
timestamp 1733704561
transform 1 0 2122 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_4
timestamp 1733704561
transform 1 0 2510 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_5
timestamp 1733704561
transform 1 0 2898 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_6
timestamp 1733704561
transform 1 0 3286 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_755577  sky130_fd_pr__pfet_01v8_lvt_755577_7
timestamp 1733704561
transform 1 0 3674 0 1 -736
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_0
timestamp 1733704561
transform 1 0 182 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_1
timestamp 1733704561
transform 1 0 552 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_2
timestamp 1733704561
transform 1 0 924 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_3
timestamp 1733704561
transform 1 0 1294 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_4
timestamp 1733704561
transform 1 0 1666 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_5
timestamp 1733704561
transform 1 0 2036 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_6
timestamp 1733704561
transform 1 0 2408 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_7
timestamp 1733704561
transform 1 0 2778 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_8
timestamp 1733704561
transform 1 0 3156 0 1 616
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_N5558H  sky130_fd_pr__pfet_01v8_lvt_N5558H_9
timestamp 1733704561
transform 1 0 3526 0 1 616
box -194 -598 194 564
use sky130_fd_pr__res_xhigh_po_0p35_5KD9UN  sky130_fd_pr__res_xhigh_po_0p35_5KD9UN_0
timestamp 1733703118
transform 1 0 4521 0 1 342
box -35 -572 35 572
use sky130_fd_pr__res_xhigh_po_0p35_5KD9UN  sky130_fd_pr__res_xhigh_po_0p35_5KD9UN_1
timestamp 1733703118
transform 1 0 4356 0 1 341
box -35 -572 35 572
<< labels >>
rlabel via2 3638 1370 3698 1430 1 VDD
port 2 n
rlabel metal2 1888 1272 1948 1332 1 i_in
port 3 n
rlabel metal2 1508 -1342 1568 -1282 1 Vinminus
port 4 n
rlabel metal2 3062 -1342 3122 -1282 1 Vinplus
port 5 n
rlabel metal2 4074 -204 4134 -144 1 Vioplus
port 6 n
rlabel metal2 4074 -100 4134 -40 1 Viominus
port 7 n
rlabel metal1 4406 1288 4466 1348 1 VSS
port 8 n
<< properties >>
string FIXED_BBOX 5468 -388 5772 928
<< end >>
