magic
tech sky130B
magscale 1 2
timestamp 1733700048
<< pwell >>
rect -296 -5773 296 5773
<< nmos >>
rect -100 4363 100 5563
rect -100 2945 100 4145
rect -100 1527 100 2727
rect -100 109 100 1309
rect -100 -1309 100 -109
rect -100 -2727 100 -1527
rect -100 -4145 100 -2945
rect -100 -5563 100 -4363
<< ndiff >>
rect -158 5551 -100 5563
rect -158 4375 -146 5551
rect -112 4375 -100 5551
rect -158 4363 -100 4375
rect 100 5551 158 5563
rect 100 4375 112 5551
rect 146 4375 158 5551
rect 100 4363 158 4375
rect -158 4133 -100 4145
rect -158 2957 -146 4133
rect -112 2957 -100 4133
rect -158 2945 -100 2957
rect 100 4133 158 4145
rect 100 2957 112 4133
rect 146 2957 158 4133
rect 100 2945 158 2957
rect -158 2715 -100 2727
rect -158 1539 -146 2715
rect -112 1539 -100 2715
rect -158 1527 -100 1539
rect 100 2715 158 2727
rect 100 1539 112 2715
rect 146 1539 158 2715
rect 100 1527 158 1539
rect -158 1297 -100 1309
rect -158 121 -146 1297
rect -112 121 -100 1297
rect -158 109 -100 121
rect 100 1297 158 1309
rect 100 121 112 1297
rect 146 121 158 1297
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1297 -146 -121
rect -112 -1297 -100 -121
rect -158 -1309 -100 -1297
rect 100 -121 158 -109
rect 100 -1297 112 -121
rect 146 -1297 158 -121
rect 100 -1309 158 -1297
rect -158 -1539 -100 -1527
rect -158 -2715 -146 -1539
rect -112 -2715 -100 -1539
rect -158 -2727 -100 -2715
rect 100 -1539 158 -1527
rect 100 -2715 112 -1539
rect 146 -2715 158 -1539
rect 100 -2727 158 -2715
rect -158 -2957 -100 -2945
rect -158 -4133 -146 -2957
rect -112 -4133 -100 -2957
rect -158 -4145 -100 -4133
rect 100 -2957 158 -2945
rect 100 -4133 112 -2957
rect 146 -4133 158 -2957
rect 100 -4145 158 -4133
rect -158 -4375 -100 -4363
rect -158 -5551 -146 -4375
rect -112 -5551 -100 -4375
rect -158 -5563 -100 -5551
rect 100 -4375 158 -4363
rect 100 -5551 112 -4375
rect 146 -5551 158 -4375
rect 100 -5563 158 -5551
<< ndiffc >>
rect -146 4375 -112 5551
rect 112 4375 146 5551
rect -146 2957 -112 4133
rect 112 2957 146 4133
rect -146 1539 -112 2715
rect 112 1539 146 2715
rect -146 121 -112 1297
rect 112 121 146 1297
rect -146 -1297 -112 -121
rect 112 -1297 146 -121
rect -146 -2715 -112 -1539
rect 112 -2715 146 -1539
rect -146 -4133 -112 -2957
rect 112 -4133 146 -2957
rect -146 -5551 -112 -4375
rect 112 -5551 146 -4375
<< psubdiff >>
rect -260 5703 -164 5737
rect 164 5703 260 5737
rect -260 5641 -226 5703
rect 226 5641 260 5703
rect -260 -5703 -226 -5641
rect 226 -5703 260 -5641
rect -260 -5737 -164 -5703
rect 164 -5737 260 -5703
<< psubdiffcont >>
rect -164 5703 164 5737
rect -260 -5641 -226 5641
rect 226 -5641 260 5641
rect -164 -5737 164 -5703
<< poly >>
rect -100 5635 100 5651
rect -100 5601 -84 5635
rect 84 5601 100 5635
rect -100 5563 100 5601
rect -100 4325 100 4363
rect -100 4291 -84 4325
rect 84 4291 100 4325
rect -100 4275 100 4291
rect -100 4217 100 4233
rect -100 4183 -84 4217
rect 84 4183 100 4217
rect -100 4145 100 4183
rect -100 2907 100 2945
rect -100 2873 -84 2907
rect 84 2873 100 2907
rect -100 2857 100 2873
rect -100 2799 100 2815
rect -100 2765 -84 2799
rect 84 2765 100 2799
rect -100 2727 100 2765
rect -100 1489 100 1527
rect -100 1455 -84 1489
rect 84 1455 100 1489
rect -100 1439 100 1455
rect -100 1381 100 1397
rect -100 1347 -84 1381
rect 84 1347 100 1381
rect -100 1309 100 1347
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1347 100 -1309
rect -100 -1381 -84 -1347
rect 84 -1381 100 -1347
rect -100 -1397 100 -1381
rect -100 -1455 100 -1439
rect -100 -1489 -84 -1455
rect 84 -1489 100 -1455
rect -100 -1527 100 -1489
rect -100 -2765 100 -2727
rect -100 -2799 -84 -2765
rect 84 -2799 100 -2765
rect -100 -2815 100 -2799
rect -100 -2873 100 -2857
rect -100 -2907 -84 -2873
rect 84 -2907 100 -2873
rect -100 -2945 100 -2907
rect -100 -4183 100 -4145
rect -100 -4217 -84 -4183
rect 84 -4217 100 -4183
rect -100 -4233 100 -4217
rect -100 -4291 100 -4275
rect -100 -4325 -84 -4291
rect 84 -4325 100 -4291
rect -100 -4363 100 -4325
rect -100 -5601 100 -5563
rect -100 -5635 -84 -5601
rect 84 -5635 100 -5601
rect -100 -5651 100 -5635
<< polycont >>
rect -84 5601 84 5635
rect -84 4291 84 4325
rect -84 4183 84 4217
rect -84 2873 84 2907
rect -84 2765 84 2799
rect -84 1455 84 1489
rect -84 1347 84 1381
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1381 84 -1347
rect -84 -1489 84 -1455
rect -84 -2799 84 -2765
rect -84 -2907 84 -2873
rect -84 -4217 84 -4183
rect -84 -4325 84 -4291
rect -84 -5635 84 -5601
<< locali >>
rect -260 5703 -164 5737
rect 164 5703 260 5737
rect -260 5641 -226 5703
rect 226 5641 260 5703
rect -100 5601 -84 5635
rect 84 5601 100 5635
rect -146 5551 -112 5567
rect -146 4359 -112 4375
rect 112 5551 146 5567
rect 112 4359 146 4375
rect -100 4291 -84 4325
rect 84 4291 100 4325
rect -100 4183 -84 4217
rect 84 4183 100 4217
rect -146 4133 -112 4149
rect -146 2941 -112 2957
rect 112 4133 146 4149
rect 112 2941 146 2957
rect -100 2873 -84 2907
rect 84 2873 100 2907
rect -100 2765 -84 2799
rect 84 2765 100 2799
rect -146 2715 -112 2731
rect -146 1523 -112 1539
rect 112 2715 146 2731
rect 112 1523 146 1539
rect -100 1455 -84 1489
rect 84 1455 100 1489
rect -100 1347 -84 1381
rect 84 1347 100 1381
rect -146 1297 -112 1313
rect -146 105 -112 121
rect 112 1297 146 1313
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1313 -112 -1297
rect 112 -121 146 -105
rect 112 -1313 146 -1297
rect -100 -1381 -84 -1347
rect 84 -1381 100 -1347
rect -100 -1489 -84 -1455
rect 84 -1489 100 -1455
rect -146 -1539 -112 -1523
rect -146 -2731 -112 -2715
rect 112 -1539 146 -1523
rect 112 -2731 146 -2715
rect -100 -2799 -84 -2765
rect 84 -2799 100 -2765
rect -100 -2907 -84 -2873
rect 84 -2907 100 -2873
rect -146 -2957 -112 -2941
rect -146 -4149 -112 -4133
rect 112 -2957 146 -2941
rect 112 -4149 146 -4133
rect -100 -4217 -84 -4183
rect 84 -4217 100 -4183
rect -100 -4325 -84 -4291
rect 84 -4325 100 -4291
rect -146 -4375 -112 -4359
rect -146 -5567 -112 -5551
rect 112 -4375 146 -4359
rect 112 -5567 146 -5551
rect -100 -5635 -84 -5601
rect 84 -5635 100 -5601
rect -260 -5703 -226 -5641
rect 226 -5703 260 -5641
rect -260 -5737 -164 -5703
rect 164 -5737 260 -5703
<< viali >>
rect -84 5601 84 5635
rect -146 4375 -112 5551
rect 112 4375 146 5551
rect -84 4291 84 4325
rect -84 4183 84 4217
rect -146 2957 -112 4133
rect 112 2957 146 4133
rect -84 2873 84 2907
rect -84 2765 84 2799
rect -146 1539 -112 2715
rect 112 1539 146 2715
rect -84 1455 84 1489
rect -84 1347 84 1381
rect -146 121 -112 1297
rect 112 121 146 1297
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1297 -112 -121
rect 112 -1297 146 -121
rect -84 -1381 84 -1347
rect -84 -1489 84 -1455
rect -146 -2715 -112 -1539
rect 112 -2715 146 -1539
rect -84 -2799 84 -2765
rect -84 -2907 84 -2873
rect -146 -4133 -112 -2957
rect 112 -4133 146 -2957
rect -84 -4217 84 -4183
rect -84 -4325 84 -4291
rect -146 -5551 -112 -4375
rect 112 -5551 146 -4375
rect -84 -5635 84 -5601
<< metal1 >>
rect -96 5635 96 5641
rect -96 5601 -84 5635
rect 84 5601 96 5635
rect -96 5595 96 5601
rect -152 5551 -106 5563
rect -152 4375 -146 5551
rect -112 4375 -106 5551
rect -152 4363 -106 4375
rect 106 5551 152 5563
rect 106 4375 112 5551
rect 146 4375 152 5551
rect 106 4363 152 4375
rect -96 4325 96 4331
rect -96 4291 -84 4325
rect 84 4291 96 4325
rect -96 4285 96 4291
rect -96 4217 96 4223
rect -96 4183 -84 4217
rect 84 4183 96 4217
rect -96 4177 96 4183
rect -152 4133 -106 4145
rect -152 2957 -146 4133
rect -112 2957 -106 4133
rect -152 2945 -106 2957
rect 106 4133 152 4145
rect 106 2957 112 4133
rect 146 2957 152 4133
rect 106 2945 152 2957
rect -96 2907 96 2913
rect -96 2873 -84 2907
rect 84 2873 96 2907
rect -96 2867 96 2873
rect -96 2799 96 2805
rect -96 2765 -84 2799
rect 84 2765 96 2799
rect -96 2759 96 2765
rect -152 2715 -106 2727
rect -152 1539 -146 2715
rect -112 1539 -106 2715
rect -152 1527 -106 1539
rect 106 2715 152 2727
rect 106 1539 112 2715
rect 146 1539 152 2715
rect 106 1527 152 1539
rect -96 1489 96 1495
rect -96 1455 -84 1489
rect 84 1455 96 1489
rect -96 1449 96 1455
rect -96 1381 96 1387
rect -96 1347 -84 1381
rect 84 1347 96 1381
rect -96 1341 96 1347
rect -152 1297 -106 1309
rect -152 121 -146 1297
rect -112 121 -106 1297
rect -152 109 -106 121
rect 106 1297 152 1309
rect 106 121 112 1297
rect 146 121 152 1297
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -1297 -146 -121
rect -112 -1297 -106 -121
rect -152 -1309 -106 -1297
rect 106 -121 152 -109
rect 106 -1297 112 -121
rect 146 -1297 152 -121
rect 106 -1309 152 -1297
rect -96 -1347 96 -1341
rect -96 -1381 -84 -1347
rect 84 -1381 96 -1347
rect -96 -1387 96 -1381
rect -96 -1455 96 -1449
rect -96 -1489 -84 -1455
rect 84 -1489 96 -1455
rect -96 -1495 96 -1489
rect -152 -1539 -106 -1527
rect -152 -2715 -146 -1539
rect -112 -2715 -106 -1539
rect -152 -2727 -106 -2715
rect 106 -1539 152 -1527
rect 106 -2715 112 -1539
rect 146 -2715 152 -1539
rect 106 -2727 152 -2715
rect -96 -2765 96 -2759
rect -96 -2799 -84 -2765
rect 84 -2799 96 -2765
rect -96 -2805 96 -2799
rect -96 -2873 96 -2867
rect -96 -2907 -84 -2873
rect 84 -2907 96 -2873
rect -96 -2913 96 -2907
rect -152 -2957 -106 -2945
rect -152 -4133 -146 -2957
rect -112 -4133 -106 -2957
rect -152 -4145 -106 -4133
rect 106 -2957 152 -2945
rect 106 -4133 112 -2957
rect 146 -4133 152 -2957
rect 106 -4145 152 -4133
rect -96 -4183 96 -4177
rect -96 -4217 -84 -4183
rect 84 -4217 96 -4183
rect -96 -4223 96 -4217
rect -96 -4291 96 -4285
rect -96 -4325 -84 -4291
rect 84 -4325 96 -4291
rect -96 -4331 96 -4325
rect -152 -4375 -106 -4363
rect -152 -5551 -146 -4375
rect -112 -5551 -106 -4375
rect -152 -5563 -106 -5551
rect 106 -4375 152 -4363
rect 106 -5551 112 -4375
rect 146 -5551 152 -4375
rect 106 -5563 152 -5551
rect -96 -5601 96 -5595
rect -96 -5635 -84 -5601
rect 84 -5635 96 -5601
rect -96 -5641 96 -5635
<< properties >>
string FIXED_BBOX -243 -5720 243 5720
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
