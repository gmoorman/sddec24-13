magic
tech sky130B
magscale 1 2
timestamp 1733686585
<< nwell >>
rect -194 -564 194 598
<< pmos >>
rect -100 -464 100 536
<< pdiff >>
rect -158 524 -100 536
rect -158 -452 -146 524
rect -112 -452 -100 524
rect -158 -464 -100 -452
rect 100 524 158 536
rect 100 -452 112 524
rect 146 -452 158 524
rect 100 -464 158 -452
<< pdiffc >>
rect -146 -452 -112 524
rect 112 -452 146 524
<< poly >>
rect -100 536 100 562
rect -100 -511 100 -464
rect -100 -545 -84 -511
rect 84 -545 100 -511
rect -100 -561 100 -545
<< polycont >>
rect -84 -545 84 -511
<< locali >>
rect -146 524 -112 540
rect -146 -468 -112 -452
rect 112 524 146 540
rect 112 -468 146 -452
rect -100 -545 -84 -511
rect 84 -545 100 -511
<< viali >>
rect -146 -452 -112 524
rect 112 -452 146 524
rect -84 -545 84 -511
<< metal1 >>
rect -152 524 -106 536
rect -152 -452 -146 524
rect -112 -452 -106 524
rect -152 -464 -106 -452
rect 106 524 152 536
rect 106 -452 112 524
rect 146 -452 152 524
rect 106 -464 152 -452
rect -96 -511 96 -505
rect -96 -545 -84 -511
rect 84 -545 96 -511
rect -96 -551 96 -545
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
