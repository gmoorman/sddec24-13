** sch_path: /home/jaxie963/caravel_pls_man_analog/caravel_user_project_analog/xschem/combination_test_DUMMY.sch
.subckt combination_test_DUMMY VDD VSS CLK Voutplus Voutminus Vioplus Viominus
*.PININFO VDD:B VSS:B CLK:B Voutplus:B Voutminus:B Vioplus:B Viominus:B
XM1 Voutplus CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=10
XM2 Voutminus CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=10
XM3 Voutplus Voutminus VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=2
XM4 Voutminus Voutplus VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=2
XM5 Voutplus CLK net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=10
XM6 Voutminus CLK net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=10
XM7 net1 Voutminus net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=2
XM8 net3 Voutplus net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=2
XM9 net2 Vioplus VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=10
XM10 net4 Viominus VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=10
.ends
.end
