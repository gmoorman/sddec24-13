magic
tech sky130B
magscale 1 2
timestamp 1731818131
<< pwell >>
rect -366 -5370 3788 -1434
<< mvpsubdiff >>
rect -300 -1512 3722 -1500
rect -300 -1612 -126 -1512
rect 3548 -1612 3722 -1512
rect -300 -1624 3722 -1612
rect -300 -1674 -176 -1624
rect -300 -5130 -288 -1674
rect -188 -5130 -176 -1674
rect -300 -5180 -176 -5130
rect 3598 -1674 3722 -1624
rect 3598 -5130 3610 -1674
rect 3710 -5130 3722 -1674
rect 3598 -5180 3722 -5130
rect -300 -5192 3722 -5180
rect -300 -5292 -126 -5192
rect 3548 -5292 3722 -5192
rect -300 -5304 3722 -5292
<< mvpsubdiffcont >>
rect -126 -1612 3548 -1512
rect -288 -5130 -188 -1674
rect 3610 -5130 3710 -1674
rect -126 -5292 3548 -5192
<< locali >>
rect -288 -1674 -188 -1512
rect -288 -5292 -188 -5130
rect 3610 -1674 3710 -1512
rect 3610 -5292 3710 -5130
<< viali >>
rect -188 -1612 -126 -1512
rect -126 -1612 3548 -1512
rect 3548 -1612 3610 -1512
rect -288 -5013 -188 -1791
rect 3610 -5013 3710 -1791
rect -188 -5292 -126 -5192
rect -126 -5292 3548 -5192
rect 3548 -5292 3610 -5192
<< metal1 >>
rect -294 -1512 3716 -1506
rect -294 -1612 -188 -1512
rect 3610 -1612 3716 -1512
rect -294 -1618 3716 -1612
rect -294 -1791 -182 -1618
rect 308 -1752 408 -1652
rect -294 -5013 -288 -1791
rect -188 -5013 -182 -1791
rect 330 -1912 382 -1752
rect 3604 -1791 3716 -1618
rect 330 -1974 382 -1964
rect 610 -1912 662 -1902
rect 610 -1974 662 -1964
rect 1450 -1912 1502 -1902
rect 1450 -1974 1502 -1964
rect 1730 -1912 1782 -1902
rect 1730 -1974 1782 -1964
rect 2570 -1912 2622 -1902
rect 2570 -1974 2622 -1964
rect 2850 -1912 2902 -1902
rect 2850 -1974 2902 -1964
rect 178 -2012 230 -2002
rect 178 -2074 230 -2064
rect 186 -2360 222 -2074
rect 254 -2112 306 -2102
rect 254 -2174 306 -2164
rect 262 -2228 298 -2174
rect 338 -2360 374 -1974
rect 458 -2012 510 -2002
rect 458 -2074 510 -2064
rect 466 -2360 502 -2074
rect 534 -2112 586 -2102
rect 534 -2174 586 -2164
rect 542 -2228 578 -2174
rect 618 -2360 654 -1974
rect 1298 -2012 1350 -2002
rect 1298 -2074 1350 -2064
rect 814 -2112 866 -2102
rect 814 -2174 866 -2164
rect 1094 -2112 1146 -2102
rect 1094 -2174 1146 -2164
rect 822 -2228 858 -2174
rect 1102 -2228 1138 -2174
rect 1306 -2360 1342 -2074
rect 1374 -2112 1426 -2102
rect 1374 -2174 1426 -2164
rect 1382 -2228 1418 -2174
rect 1458 -2360 1494 -1974
rect 1578 -2012 1630 -2002
rect 1578 -2074 1630 -2064
rect 1586 -2360 1622 -2074
rect 1654 -2112 1706 -2102
rect 1654 -2174 1706 -2164
rect 1662 -2228 1698 -2174
rect 1738 -2360 1774 -1974
rect 2418 -2012 2470 -2002
rect 2418 -2074 2470 -2064
rect 1934 -2112 1986 -2102
rect 1934 -2174 1986 -2164
rect 2214 -2112 2266 -2102
rect 2214 -2174 2266 -2164
rect 1942 -2228 1978 -2174
rect 2222 -2228 2258 -2174
rect 2426 -2360 2462 -2074
rect 2494 -2112 2546 -2102
rect 2494 -2174 2546 -2164
rect 2502 -2228 2538 -2174
rect 2578 -2360 2614 -1974
rect 2698 -2012 2750 -2002
rect 2698 -2074 2750 -2064
rect 2706 -2360 2742 -2074
rect 2774 -2112 2826 -2102
rect 2774 -2174 2826 -2164
rect 2782 -2228 2818 -2174
rect 2858 -2360 2894 -1974
rect 3220 -2010 3320 -1978
rect 2960 -2062 2970 -2010
rect 3022 -2062 3320 -2010
rect 3220 -2078 3320 -2062
rect 262 -2798 298 -2738
rect 542 -2798 578 -2738
rect 746 -2822 782 -2640
rect 822 -2798 858 -2738
rect 178 -2836 230 -2826
rect 178 -2898 230 -2888
rect 458 -2836 510 -2826
rect 458 -2898 510 -2888
rect 738 -2832 790 -2822
rect 738 -2894 790 -2884
rect 186 -4298 222 -2898
rect 330 -2936 382 -2926
rect 330 -2998 382 -2988
rect 262 -3082 298 -3022
rect 338 -3180 374 -2998
rect 466 -3180 502 -2898
rect 898 -2926 934 -2640
rect 1026 -2822 1062 -2640
rect 1102 -2798 1138 -2738
rect 1018 -2832 1070 -2822
rect 1018 -2894 1070 -2884
rect 1178 -2926 1214 -2640
rect 1382 -2798 1418 -2738
rect 1662 -2798 1698 -2738
rect 1866 -2822 1902 -2640
rect 1942 -2798 1978 -2738
rect 1298 -2836 1350 -2826
rect 1298 -2898 1350 -2888
rect 1578 -2836 1630 -2826
rect 1578 -2898 1630 -2888
rect 1858 -2832 1910 -2822
rect 1858 -2894 1910 -2884
rect 610 -2936 662 -2926
rect 610 -2998 662 -2988
rect 890 -2936 942 -2926
rect 890 -2998 942 -2988
rect 1170 -2936 1222 -2926
rect 1170 -2998 1222 -2988
rect 542 -3082 578 -3022
rect 618 -3180 654 -2998
rect 822 -3082 858 -3022
rect 1102 -3082 1138 -3022
rect 1306 -3180 1342 -2898
rect 1450 -2936 1502 -2926
rect 1450 -2998 1502 -2988
rect 1382 -3082 1418 -3022
rect 1458 -3180 1494 -2998
rect 1586 -3180 1622 -2898
rect 2018 -2926 2054 -2640
rect 2146 -2822 2182 -2640
rect 2222 -2798 2258 -2738
rect 2138 -2832 2190 -2822
rect 2138 -2894 2190 -2884
rect 2298 -2926 2334 -2640
rect 2502 -2798 2538 -2738
rect 2782 -2798 2818 -2738
rect 2418 -2836 2470 -2826
rect 2418 -2898 2470 -2888
rect 2698 -2836 2750 -2826
rect 3198 -2838 3298 -2812
rect 2698 -2898 2750 -2888
rect 2850 -2890 3298 -2838
rect 1730 -2936 1782 -2926
rect 1730 -2998 1782 -2988
rect 2010 -2936 2062 -2926
rect 2010 -2998 2062 -2988
rect 2290 -2936 2342 -2926
rect 2290 -2998 2342 -2988
rect 1662 -3082 1698 -3022
rect 1738 -3180 1774 -2998
rect 1942 -3082 1978 -3022
rect 2222 -3082 2258 -3022
rect 2426 -3180 2462 -2898
rect 2570 -2936 2622 -2926
rect 2570 -2998 2622 -2988
rect 2502 -3082 2538 -3022
rect 2578 -3180 2614 -2998
rect 2706 -3180 2742 -2898
rect 2850 -2936 2902 -2890
rect 3198 -2912 3298 -2890
rect 2850 -2998 2902 -2988
rect 2782 -3082 2818 -3022
rect 2858 -3180 2894 -2998
rect 262 -3646 298 -3592
rect 542 -3646 578 -3592
rect 254 -3656 306 -3646
rect 254 -3718 306 -3708
rect 534 -3656 586 -3646
rect 534 -3718 586 -3708
rect 746 -3846 782 -3460
rect 822 -3646 858 -3592
rect 814 -3656 866 -3646
rect 814 -3718 866 -3708
rect 898 -3746 934 -3460
rect 890 -3756 942 -3746
rect 890 -3818 942 -3808
rect 1026 -3846 1062 -3460
rect 1102 -3646 1138 -3592
rect 1094 -3656 1146 -3646
rect 1094 -3718 1146 -3708
rect 1178 -3746 1214 -3460
rect 1382 -3646 1418 -3592
rect 1662 -3646 1698 -3592
rect 1374 -3656 1426 -3646
rect 1374 -3718 1426 -3708
rect 1654 -3656 1706 -3646
rect 1654 -3718 1706 -3708
rect 1170 -3756 1222 -3746
rect 1170 -3818 1222 -3808
rect 1866 -3846 1902 -3460
rect 1942 -3646 1978 -3592
rect 1934 -3656 1986 -3646
rect 1934 -3718 1986 -3708
rect 2018 -3746 2054 -3460
rect 2010 -3756 2062 -3746
rect 2010 -3818 2062 -3808
rect 2146 -3846 2182 -3460
rect 2222 -3646 2258 -3592
rect 2214 -3656 2266 -3646
rect 2214 -3718 2266 -3708
rect 2298 -3746 2334 -3460
rect 2502 -3646 2538 -3592
rect 2782 -3646 2818 -3592
rect 2494 -3656 2546 -3646
rect 2494 -3718 2546 -3708
rect 2774 -3656 2826 -3646
rect 2774 -3718 2826 -3708
rect 2290 -3756 2342 -3746
rect 2290 -3818 2342 -3808
rect 738 -3856 790 -3846
rect 738 -4244 790 -3908
rect 1018 -3856 1070 -3846
rect 1018 -3918 1070 -3908
rect 1858 -3856 1910 -3846
rect 1858 -3918 1910 -3908
rect 2138 -3856 2190 -3846
rect 2138 -3918 2190 -3908
rect 154 -4398 254 -4298
rect 714 -4344 814 -4244
rect -294 -5186 -182 -5013
rect 418 -5186 428 -4886
rect 906 -4994 1006 -4894
rect 928 -5186 982 -4994
rect 2994 -5186 3004 -4886
rect 3604 -5013 3610 -1791
rect 3710 -5013 3716 -1791
rect 3604 -5186 3716 -5013
rect -294 -5192 3716 -5186
rect -294 -5292 -188 -5192
rect 3610 -5292 3716 -5192
rect -294 -5298 3716 -5292
<< via1 >>
rect 330 -1964 382 -1912
rect 610 -1964 662 -1912
rect 1450 -1964 1502 -1912
rect 1730 -1964 1782 -1912
rect 2570 -1964 2622 -1912
rect 2850 -1964 2902 -1912
rect 178 -2064 230 -2012
rect 254 -2164 306 -2112
rect 458 -2064 510 -2012
rect 534 -2164 586 -2112
rect 1298 -2064 1350 -2012
rect 814 -2164 866 -2112
rect 1094 -2164 1146 -2112
rect 1374 -2164 1426 -2112
rect 1578 -2064 1630 -2012
rect 1654 -2164 1706 -2112
rect 2418 -2064 2470 -2012
rect 1934 -2164 1986 -2112
rect 2214 -2164 2266 -2112
rect 2494 -2164 2546 -2112
rect 2698 -2064 2750 -2012
rect 2774 -2164 2826 -2112
rect 2970 -2062 3022 -2010
rect 178 -2888 230 -2836
rect 458 -2888 510 -2836
rect 738 -2884 790 -2832
rect 330 -2988 382 -2936
rect 1018 -2884 1070 -2832
rect 1298 -2888 1350 -2836
rect 1578 -2888 1630 -2836
rect 1858 -2884 1910 -2832
rect 610 -2988 662 -2936
rect 890 -2988 942 -2936
rect 1170 -2988 1222 -2936
rect 1450 -2988 1502 -2936
rect 2138 -2884 2190 -2832
rect 2418 -2888 2470 -2836
rect 2698 -2888 2750 -2836
rect 1730 -2988 1782 -2936
rect 2010 -2988 2062 -2936
rect 2290 -2988 2342 -2936
rect 2570 -2988 2622 -2936
rect 2850 -2988 2902 -2936
rect 254 -3708 306 -3656
rect 534 -3708 586 -3656
rect 814 -3708 866 -3656
rect 890 -3808 942 -3756
rect 1094 -3708 1146 -3656
rect 1374 -3708 1426 -3656
rect 1654 -3708 1706 -3656
rect 1170 -3808 1222 -3756
rect 1934 -3708 1986 -3656
rect 2010 -3808 2062 -3756
rect 2214 -3708 2266 -3656
rect 2494 -3708 2546 -3656
rect 2774 -3708 2826 -3656
rect 2290 -3808 2342 -3756
rect 738 -3908 790 -3856
rect 1018 -3908 1070 -3856
rect 1858 -3908 1910 -3856
rect 2138 -3908 2190 -3856
rect -182 -5186 418 -4886
rect 3004 -5186 3604 -4886
<< metal2 >>
rect 320 -1964 330 -1912
rect 382 -1964 610 -1912
rect 662 -1964 1450 -1912
rect 1502 -1964 1730 -1912
rect 1782 -1964 2570 -1912
rect 2622 -1964 2850 -1912
rect 2902 -1964 3104 -1912
rect 2970 -2010 3022 -2000
rect -76 -2064 178 -2012
rect 230 -2064 458 -2012
rect 510 -2064 1298 -2012
rect 1350 -2064 1578 -2012
rect 1630 -2064 2418 -2012
rect 2470 -2064 2698 -2012
rect 2750 -2064 2760 -2012
rect -76 -3856 -24 -2064
rect 2970 -2112 3022 -2062
rect 58 -2164 254 -2112
rect 306 -2164 534 -2112
rect 586 -2164 814 -2112
rect 866 -2164 1094 -2112
rect 1146 -2164 1374 -2112
rect 1426 -2164 1654 -2112
rect 1706 -2164 1934 -2112
rect 1986 -2164 2214 -2112
rect 2266 -2164 2494 -2112
rect 2546 -2164 2774 -2112
rect 2826 -2164 3022 -2112
rect 58 -3656 110 -2164
rect 728 -2836 738 -2832
rect 168 -2888 178 -2836
rect 230 -2888 458 -2836
rect 510 -2884 738 -2836
rect 790 -2836 800 -2832
rect 1008 -2836 1018 -2832
rect 790 -2884 1018 -2836
rect 1070 -2836 1080 -2832
rect 1848 -2836 1858 -2832
rect 1070 -2884 1298 -2836
rect 510 -2888 1298 -2884
rect 1350 -2888 1578 -2836
rect 1630 -2884 1858 -2836
rect 1910 -2836 1920 -2832
rect 2128 -2836 2138 -2832
rect 1910 -2884 2138 -2836
rect 2190 -2836 2200 -2832
rect 2190 -2884 2418 -2836
rect 1630 -2888 2418 -2884
rect 2470 -2888 2698 -2836
rect 2750 -2888 2760 -2836
rect 320 -2988 330 -2936
rect 382 -2988 610 -2936
rect 662 -2988 890 -2936
rect 942 -2988 1170 -2936
rect 1222 -2988 1450 -2936
rect 1502 -2988 1730 -2936
rect 1782 -2988 2010 -2936
rect 2062 -2988 2290 -2936
rect 2342 -2988 2570 -2936
rect 2622 -2988 2850 -2936
rect 2902 -2988 2912 -2936
rect 330 -2990 2902 -2988
rect 2970 -3656 3022 -2164
rect 58 -3708 254 -3656
rect 306 -3708 534 -3656
rect 586 -3708 814 -3656
rect 866 -3708 1094 -3656
rect 1146 -3708 1374 -3656
rect 1426 -3708 1654 -3656
rect 1706 -3708 1934 -3656
rect 1986 -3708 2214 -3656
rect 2266 -3708 2494 -3656
rect 2546 -3708 2774 -3656
rect 2826 -3708 3022 -3656
rect 3052 -3756 3104 -1964
rect 880 -3808 890 -3756
rect 942 -3808 1170 -3756
rect 1222 -3808 2010 -3756
rect 2062 -3808 2290 -3756
rect 2342 -3808 3104 -3756
rect -76 -3908 738 -3856
rect 790 -3908 1018 -3856
rect 1070 -3908 1858 -3856
rect 1910 -3908 2138 -3856
rect 2190 -3908 2200 -3856
rect -182 -4886 418 -4876
rect -182 -5196 418 -5186
rect 3004 -4886 3604 -4876
rect 3004 -5196 3604 -5186
<< via2 >>
rect -182 -5186 418 -4886
rect 3004 -5186 3604 -4886
<< metal3 >>
rect -192 -4886 428 -4881
rect -192 -5186 -182 -4886
rect 418 -5186 428 -4886
rect -192 -5191 428 -5186
rect 2994 -4886 3614 -4881
rect 2994 -5186 3004 -4886
rect 3604 -5186 3614 -4886
rect 2994 -5191 3614 -5186
<< via3 >>
rect -182 -5186 418 -4886
rect 3004 -5186 3604 -4886
<< metal4 >>
rect -183 -4886 419 -4885
rect -183 -5186 -182 -4886
rect 418 -5186 419 -4886
rect -183 -5187 419 -5186
rect 3003 -4886 3605 -4885
rect 3003 -5186 3004 -4886
rect 3604 -5186 3605 -4886
rect 3003 -5187 3605 -5186
use sky130_fd_pr__nfet_01v8_PHZV97  xm25
timestamp 1731817339
transform 1 0 280 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm26
timestamp 1731817339
transform 1 0 560 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm27
timestamp 1731817339
transform 1 0 840 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm28
timestamp 1731817339
transform 1 0 1120 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm29
timestamp 1731817339
transform 1 0 1400 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm30
timestamp 1731817339
transform 1 0 1680 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm31
timestamp 1731817339
transform 1 0 1960 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm32
timestamp 1731817339
transform 1 0 2240 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm33
timestamp 1731817339
transform 1 0 2520 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm34
timestamp 1731817339
transform 1 0 2800 0 1 -2500
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm35
timestamp 1731817339
transform 1 0 280 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm36
timestamp 1731817339
transform 1 0 560 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm37
timestamp 1731817339
transform 1 0 840 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm38
timestamp 1731817339
transform 1 0 1120 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm39
timestamp 1731817339
transform 1 0 1400 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm40
timestamp 1731817339
transform 1 0 1680 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm41
timestamp 1731817339
transform 1 0 1960 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm42
timestamp 1731817339
transform 1 0 2240 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm43
timestamp 1731817339
transform 1 0 2520 0 1 -3320
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm44
timestamp 1731817339
transform 1 0 2800 0 1 -3320
box -73 -288 73 288
<< labels >>
rlabel metal1 154 -4398 254 -4298 1 M7_net
port 1 n
rlabel metal1 714 -4344 814 -4244 1 M8_net
port 2 n
rlabel metal1 3198 -2912 3298 -2812 1 voutplus
port 3 n
rlabel metal1 308 -1752 408 -1652 1 voutminus
port 4 n
rlabel metal1 3220 -2078 3320 -1978 1 CLK
port 5 n
rlabel metal1 906 -4994 1006 -4894 1 VSS
port 6 n
<< properties >>
string FIXED_BBOX -238 -5242 3660 -1562
<< end >>
