magic
tech sky130B
magscale 1 2
timestamp 1726587868
<< pwell >>
rect -140 680 416 2596
<< mvnmos >>
rect 88 938 188 2338
<< mvndiff >>
rect 30 2326 88 2338
rect 30 950 42 2326
rect 76 950 88 2326
rect 30 938 88 950
rect 188 2326 246 2338
rect 188 950 200 2326
rect 234 950 246 2326
rect 188 938 246 950
<< mvndiffc >>
rect 42 950 76 2326
rect 200 950 234 2326
<< mvpsubdiff >>
rect -104 2548 380 2560
rect -104 2514 4 2548
rect 272 2514 380 2548
rect -104 2502 380 2514
rect -104 2452 -46 2502
rect -104 824 -92 2452
rect -58 824 -46 2452
rect 322 2452 380 2502
rect -104 774 -46 824
rect 322 824 334 2452
rect 368 824 380 2452
rect 322 774 380 824
rect -104 762 380 774
rect -104 728 4 762
rect 272 728 380 762
rect -104 716 380 728
<< mvpsubdiffcont >>
rect 4 2514 272 2548
rect -92 824 -58 2452
rect 334 824 368 2452
rect 4 728 272 762
<< poly >>
rect 88 2410 188 2426
rect 88 2376 104 2410
rect 172 2376 188 2410
rect 88 2338 188 2376
rect 88 900 188 938
rect 88 866 104 900
rect 172 866 188 900
rect 88 850 188 866
<< polycont >>
rect 104 2376 172 2410
rect 104 866 172 900
<< locali >>
rect -100 2548 380 2560
rect -100 2514 4 2548
rect 272 2514 380 2548
rect -100 2500 380 2514
rect -100 2452 -40 2500
rect -100 824 -92 2452
rect -58 824 -40 2452
rect 320 2452 380 2500
rect 88 2376 104 2410
rect 172 2376 188 2410
rect 42 2326 76 2342
rect 42 934 76 950
rect 200 2326 234 2342
rect 200 934 234 950
rect 88 866 104 900
rect 172 866 188 900
rect -100 762 -40 824
rect 320 824 334 2452
rect 368 824 380 2452
rect 320 762 380 824
rect -100 728 4 762
rect 272 728 380 762
rect -100 680 380 728
rect -100 480 180 680
rect 340 480 380 680
rect -100 420 380 480
<< viali >>
rect 104 2376 172 2410
rect 42 950 76 2326
rect 200 950 234 2326
rect 104 866 172 900
rect 180 480 340 680
<< metal1 >>
rect 120 2416 160 2420
rect 92 2410 184 2416
rect 92 2376 104 2410
rect 172 2376 184 2410
rect 92 2370 184 2376
rect 36 2326 82 2338
rect 36 1896 42 2326
rect -24 1832 -14 1896
rect 36 950 42 1832
rect 76 950 82 2326
rect 36 938 82 950
rect 120 906 160 2370
rect 194 2326 240 2338
rect 194 950 200 2326
rect 234 1760 240 2326
rect 234 1520 440 1760
rect 234 950 240 1520
rect 194 938 240 950
rect 92 900 184 906
rect 90 840 100 900
rect 180 840 190 900
rect -100 680 380 740
rect -100 480 180 680
rect 340 480 380 680
rect -100 420 380 480
<< via1 >>
rect -14 1832 42 1896
rect 42 1832 72 1896
rect 100 866 104 900
rect 104 866 172 900
rect 172 866 180 900
rect 100 840 180 866
<< reram >>
rect 226 1546 426 1746
<< metal2 >>
rect -80 2820 120 2830
rect -80 2610 120 2620
rect -20 1906 60 2610
rect -20 1896 72 1906
rect -20 1840 -14 1896
rect -14 1822 72 1832
rect 200 1746 440 1760
rect 200 1546 226 1746
rect 426 1680 440 1746
rect 580 1740 780 1750
rect 426 1600 580 1680
rect 426 1546 440 1600
rect 200 1520 440 1546
rect 580 1530 780 1540
rect -360 900 -160 960
rect 100 900 180 910
rect -360 840 100 900
rect -360 760 -160 840
rect 100 830 180 840
<< via2 >>
rect -80 2620 120 2820
rect 580 1540 780 1740
<< metal3 >>
rect -90 2820 130 2825
rect -90 2620 -80 2820
rect 120 2620 130 2820
rect -90 2615 130 2620
rect 570 1740 790 1745
rect 570 1540 580 1740
rect 780 1540 790 1740
rect 570 1535 790 1540
<< labels >>
flabel metal1 -60 480 140 680 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal2 -360 760 -160 960 0 FreeSans 256 0 0 0 WL
port 2 nsew
flabel metal3 580 1540 780 1740 0 FreeSans 256 0 0 0 BL
port 3 nsew
flabel metal3 -80 2620 120 2820 0 FreeSans 256 0 0 0 SL
port 0 nsew
flabel metal1 226 1546 426 1746 0 FreeSans 256 0 0 0 XR1.BE
flabel reram 226 1546 426 1746 0 FreeSans 256 0 0 0 XR1.TE
<< end >>
