magic
tech sky130B
magscale 1 2
timestamp 1733718626
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 2 67 813 203
rect 29 21 813 67
rect 29 -17 63 21
<< scnmos >>
rect 80 93 110 177
rect 281 47 311 177
rect 365 47 395 177
rect 449 47 479 177
rect 533 47 563 177
rect 617 47 647 177
rect 701 47 731 177
<< scpmoshvt >>
rect 80 297 110 381
rect 177 297 207 497
rect 261 297 291 497
rect 449 297 479 497
rect 533 297 563 497
rect 617 297 647 497
rect 701 297 731 497
<< ndiff >>
rect 28 149 80 177
rect 28 115 36 149
rect 70 115 80 149
rect 28 93 80 115
rect 110 149 162 177
rect 110 115 120 149
rect 154 115 162 149
rect 110 93 162 115
rect 229 163 281 177
rect 229 129 237 163
rect 271 129 281 163
rect 229 95 281 129
rect 229 61 237 95
rect 271 61 281 95
rect 229 47 281 61
rect 311 163 365 177
rect 311 129 321 163
rect 355 129 365 163
rect 311 47 365 129
rect 395 163 449 177
rect 395 129 405 163
rect 439 129 449 163
rect 395 95 449 129
rect 395 61 405 95
rect 439 61 449 95
rect 395 47 449 61
rect 479 95 533 177
rect 479 61 489 95
rect 523 61 533 95
rect 479 47 533 61
rect 563 163 617 177
rect 563 129 573 163
rect 607 129 617 163
rect 563 95 617 129
rect 563 61 573 95
rect 607 61 617 95
rect 563 47 617 61
rect 647 95 701 177
rect 647 61 657 95
rect 691 61 701 95
rect 647 47 701 61
rect 731 163 787 177
rect 731 129 741 163
rect 775 129 787 163
rect 731 95 787 129
rect 731 61 741 95
rect 775 61 787 95
rect 731 47 787 61
<< pdiff >>
rect 125 477 177 497
rect 125 443 133 477
rect 167 443 177 477
rect 125 409 177 443
rect 125 381 133 409
rect 28 362 80 381
rect 28 328 36 362
rect 70 328 80 362
rect 28 297 80 328
rect 110 375 133 381
rect 167 375 177 409
rect 110 297 177 375
rect 207 477 261 497
rect 207 443 217 477
rect 251 443 261 477
rect 207 409 261 443
rect 207 375 217 409
rect 251 375 261 409
rect 207 341 261 375
rect 207 307 217 341
rect 251 307 261 341
rect 207 297 261 307
rect 291 477 343 497
rect 291 443 301 477
rect 335 443 343 477
rect 291 409 343 443
rect 291 375 301 409
rect 335 375 343 409
rect 291 297 343 375
rect 397 477 449 497
rect 397 443 405 477
rect 439 443 449 477
rect 397 409 449 443
rect 397 375 405 409
rect 439 375 449 409
rect 397 297 449 375
rect 479 409 533 497
rect 479 375 489 409
rect 523 375 533 409
rect 479 341 533 375
rect 479 307 489 341
rect 523 307 533 341
rect 479 297 533 307
rect 563 477 617 497
rect 563 443 573 477
rect 607 443 617 477
rect 563 409 617 443
rect 563 375 573 409
rect 607 375 617 409
rect 563 341 617 375
rect 563 307 573 341
rect 607 307 617 341
rect 563 297 617 307
rect 647 485 701 497
rect 647 451 657 485
rect 691 451 701 485
rect 647 417 701 451
rect 647 383 657 417
rect 691 383 701 417
rect 647 297 701 383
rect 731 477 787 497
rect 731 443 741 477
rect 775 443 787 477
rect 731 409 787 443
rect 731 375 741 409
rect 775 375 787 409
rect 731 341 787 375
rect 731 307 741 341
rect 775 307 787 341
rect 731 297 787 307
<< ndiffc >>
rect 36 115 70 149
rect 120 115 154 149
rect 237 129 271 163
rect 237 61 271 95
rect 321 129 355 163
rect 405 129 439 163
rect 405 61 439 95
rect 489 61 523 95
rect 573 129 607 163
rect 573 61 607 95
rect 657 61 691 95
rect 741 129 775 163
rect 741 61 775 95
<< pdiffc >>
rect 133 443 167 477
rect 36 328 70 362
rect 133 375 167 409
rect 217 443 251 477
rect 217 375 251 409
rect 217 307 251 341
rect 301 443 335 477
rect 301 375 335 409
rect 405 443 439 477
rect 405 375 439 409
rect 489 375 523 409
rect 489 307 523 341
rect 573 443 607 477
rect 573 375 607 409
rect 573 307 607 341
rect 657 451 691 485
rect 657 383 691 417
rect 741 443 775 477
rect 741 375 775 409
rect 741 307 775 341
<< poly >>
rect 177 497 207 523
rect 261 497 291 523
rect 449 497 479 523
rect 533 497 563 523
rect 617 497 647 523
rect 701 497 731 523
rect 80 381 110 407
rect 80 265 110 297
rect 35 249 110 265
rect 35 215 54 249
rect 88 215 110 249
rect 35 199 110 215
rect 177 265 207 297
rect 261 265 291 297
rect 449 265 479 297
rect 533 265 563 297
rect 177 249 395 265
rect 177 215 217 249
rect 251 215 395 249
rect 177 199 395 215
rect 80 177 110 199
rect 281 177 311 199
rect 365 177 395 199
rect 449 249 563 265
rect 449 215 489 249
rect 523 215 563 249
rect 449 199 563 215
rect 449 177 479 199
rect 533 177 563 199
rect 617 265 647 297
rect 701 265 731 297
rect 617 249 731 265
rect 617 215 668 249
rect 702 215 731 249
rect 617 199 731 215
rect 617 177 647 199
rect 701 177 731 199
rect 80 67 110 93
rect 281 21 311 47
rect 365 21 395 47
rect 449 21 479 47
rect 533 21 563 47
rect 617 21 647 47
rect 701 21 731 47
<< polycont >>
rect 54 215 88 249
rect 217 215 251 249
rect 489 215 523 249
rect 668 215 702 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 117 477 183 527
rect 117 443 133 477
rect 167 443 183 477
rect 117 409 183 443
rect 36 362 70 383
rect 117 375 133 409
rect 167 375 183 409
rect 217 477 251 493
rect 217 409 251 443
rect 217 341 251 375
rect 294 477 344 527
rect 294 443 301 477
rect 335 443 344 477
rect 294 409 344 443
rect 294 375 301 409
rect 335 375 344 409
rect 294 359 344 375
rect 391 477 607 493
rect 391 443 405 477
rect 439 459 573 477
rect 439 443 447 459
rect 391 409 447 443
rect 391 375 405 409
rect 439 375 447 409
rect 391 359 447 375
rect 481 409 530 425
rect 481 375 489 409
rect 523 375 530 409
rect 70 328 173 333
rect 36 299 173 328
rect 17 249 105 265
rect 17 215 54 249
rect 88 215 105 249
rect 17 199 105 215
rect 139 249 173 299
rect 481 341 530 375
rect 481 323 489 341
rect 251 307 489 323
rect 523 307 530 341
rect 217 289 530 307
rect 573 409 607 443
rect 573 341 607 375
rect 641 485 707 527
rect 641 451 657 485
rect 691 451 707 485
rect 641 417 707 451
rect 641 383 657 417
rect 691 383 707 417
rect 641 367 707 383
rect 741 477 796 493
rect 775 443 796 477
rect 741 409 796 443
rect 775 375 796 409
rect 741 341 796 375
rect 607 307 741 333
rect 775 307 796 341
rect 573 291 796 307
rect 139 215 217 249
rect 251 215 267 249
rect 139 165 173 215
rect 305 181 356 289
rect 390 249 618 255
rect 390 215 489 249
rect 523 215 618 249
rect 652 249 811 255
rect 652 215 668 249
rect 702 215 811 249
rect 36 149 70 165
rect 36 17 70 115
rect 120 149 173 165
rect 154 115 173 149
rect 120 89 173 115
rect 215 163 271 181
rect 215 129 237 163
rect 305 163 371 181
rect 305 129 321 163
rect 355 129 371 163
rect 405 163 796 181
rect 439 145 573 163
rect 439 129 455 145
rect 215 95 271 129
rect 405 95 455 129
rect 557 129 573 145
rect 607 145 741 163
rect 607 129 623 145
rect 215 61 237 95
rect 271 61 405 95
rect 439 61 455 95
rect 215 51 455 61
rect 489 95 523 111
rect 489 17 523 61
rect 557 95 623 129
rect 725 129 741 145
rect 775 129 796 163
rect 557 61 573 95
rect 607 61 623 95
rect 557 51 623 61
rect 657 95 691 111
rect 657 17 691 61
rect 725 95 796 129
rect 725 61 741 95
rect 775 61 796 95
rect 725 53 796 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 B1_N
port 6 nsew
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel locali s 489 221 523 255 0 FreeSans 400 180 0 0 A2
port 8 nsew
flabel locali s 673 221 707 255 0 FreeSans 400 180 0 0 A1
port 9 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 o21bai_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string path 0.000 0.000 4.140 0.000 
<< end >>
