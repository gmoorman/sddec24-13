magic
tech sky130B
magscale 1 2
timestamp 1733715975
<< nwell >>
rect -999 10715 3920 16360
<< pwell >>
rect 4931 10594 7846 13215
rect 1446 9209 7846 10594
rect 1446 9185 5167 9209
rect 1446 9154 5154 9185
rect 5157 9154 5306 9178
rect 1446 9095 5306 9154
rect 5316 9126 7846 9209
rect 1446 8654 5300 9095
rect 5310 8685 7846 9126
rect 1446 8234 5326 8654
rect 5336 8234 7846 8685
rect 1446 8066 7846 8234
<< mvpsubdiff >>
rect 5173 9131 5297 9177
rect 5173 8226 5185 9131
rect 5285 8226 5297 9131
rect 5173 8188 5297 8226
<< mvnsubdiff >>
rect -752 15642 -628 15666
rect -752 15296 -740 15642
rect -640 15296 -628 15642
rect -752 15272 -628 15296
<< mvpsubdiffcont >>
rect 5185 8226 5285 9131
<< mvnsubdiffcont >>
rect -740 15296 -640 15642
<< locali >>
rect -758 15642 -618 15675
rect -758 15296 -740 15642
rect -640 15296 -618 15642
rect -758 15268 -618 15296
rect 5185 9131 5285 9154
rect 5185 8203 5285 8226
<< viali >>
rect -740 15353 -640 15491
rect 5185 8478 5285 8879
<< metal1 >>
rect 1660 16480 1760 16500
rect 1660 16420 1680 16480
rect 1740 16420 1760 16480
rect -746 15620 -634 15666
rect -20 15620 100 16020
rect 160 15852 300 15860
rect 160 15800 200 15852
rect 252 15800 300 15852
rect 540 15852 680 15860
rect 540 15800 600 15852
rect 652 15800 680 15852
rect -1240 15520 100 15620
rect -746 15491 -634 15520
rect -746 15353 -740 15491
rect -640 15353 -634 15491
rect -746 15279 -634 15353
rect -20 13820 100 15520
rect -20 13760 20 13820
rect 80 13760 100 13820
rect -20 13740 100 13760
rect -400 13092 -280 13120
rect -400 13040 -360 13092
rect -308 13040 -280 13092
rect -800 10660 -660 11340
rect -400 11300 -280 13040
rect 360 13072 480 15740
rect 740 13820 860 16020
rect 960 16012 1040 16040
rect 960 15960 980 16012
rect 1032 15960 1042 16012
rect 960 15860 1040 15960
rect 1660 15860 1760 16420
rect 2380 16012 2460 16040
rect 2380 15960 2400 16012
rect 2452 15960 2462 16012
rect 920 15800 1060 15860
rect 1300 15852 1440 15860
rect 1300 15800 1340 15852
rect 1392 15800 1440 15852
rect 1660 15800 1680 15860
rect 1740 15800 1760 15860
rect 1960 15852 2100 15860
rect 1960 15800 2000 15852
rect 2052 15800 2100 15852
rect 2380 15800 2460 15960
rect 1100 13980 1260 15740
rect 740 13760 780 13820
rect 840 13760 860 13820
rect 740 13740 860 13760
rect 1500 13160 1620 15760
rect 1800 13420 1920 15760
rect 2160 13980 2280 15740
rect 2540 13820 2660 16020
rect 2720 15852 2860 15860
rect 2720 15800 2760 15852
rect 2812 15800 2860 15852
rect 3100 15852 3240 15860
rect 3100 15800 3140 15852
rect 3192 15800 3240 15852
rect 2540 13760 2580 13820
rect 2640 13760 2660 13820
rect 2540 13740 2660 13760
rect 2920 13640 3040 15740
rect 3300 13820 3420 16020
rect 3480 15852 3620 15860
rect 3480 15800 3520 15852
rect 3572 15800 3620 15852
rect 3300 13760 3340 13820
rect 3400 13760 3420 13820
rect 3300 13740 3420 13760
rect 2920 13580 2960 13640
rect 3020 13580 3040 13640
rect 2920 13560 3040 13580
rect 3680 13640 3800 14140
rect 3680 13580 3720 13640
rect 3780 13580 3800 13640
rect 3680 13560 3800 13580
rect 6500 13640 6600 13660
rect 6500 13580 6520 13640
rect 6580 13580 6600 13640
rect 1800 13360 1840 13420
rect 1900 13360 1920 13420
rect 1800 13340 1920 13360
rect 2260 13420 2380 13440
rect 2260 13360 2300 13420
rect 2360 13360 2380 13420
rect 360 13020 400 13072
rect 452 13020 480 13072
rect -580 11092 -480 11240
rect -580 11040 -560 11092
rect -508 11040 -480 11092
rect -580 11020 -480 11040
rect -380 11080 -280 11100
rect -380 11020 -360 11080
rect -300 11020 -280 11080
rect -200 11092 -100 11240
rect -200 11040 -180 11092
rect -128 11040 -100 11092
rect -200 11020 -100 11040
rect -800 10600 -760 10660
rect -700 10600 -660 10660
rect -800 10580 -660 10600
rect -380 10440 -280 11020
rect -20 10660 100 12860
rect 360 11300 480 13020
rect 1120 13072 1240 13120
rect 1500 13100 1540 13160
rect 1600 13100 1620 13160
rect 1500 13080 1620 13100
rect 1877 13160 2004 13183
rect 1877 13100 1920 13160
rect 1980 13100 2004 13160
rect 1120 13020 1160 13072
rect 1212 13020 1240 13072
rect 180 11092 280 11240
rect 180 11040 200 11092
rect 252 11040 280 11092
rect 180 11020 280 11040
rect 560 11092 660 11220
rect 560 11040 580 11092
rect 632 11040 660 11092
rect 560 11020 660 11040
rect 740 10840 860 12860
rect 1120 11300 1240 13020
rect 940 11092 1040 11220
rect 940 11040 960 11092
rect 1012 11040 1040 11092
rect 940 11020 1040 11040
rect 1160 11080 1280 11100
rect 1160 11020 1180 11080
rect 1240 11020 1280 11080
rect 1320 11092 1420 11220
rect 1320 11040 1340 11092
rect 1392 11040 1420 11092
rect 1320 11020 1420 11040
rect 740 10780 780 10840
rect 840 10780 860 10840
rect 740 10760 860 10780
rect -20 10600 0 10660
rect 60 10600 100 10660
rect -20 10580 100 10600
rect -380 10380 -360 10440
rect -300 10380 -280 10440
rect -380 10360 -280 10380
rect 1160 10280 1280 11020
rect 1160 10220 1180 10280
rect 1240 10220 1280 10280
rect 1160 10200 1280 10220
rect 1500 10840 1620 11420
rect 1877 11097 2004 13100
rect 2260 11140 2380 13360
rect 5240 13400 5380 13440
rect 5240 13340 5280 13400
rect 5340 13340 5380 13400
rect 5240 13260 5380 13340
rect 5880 13420 6000 13440
rect 5880 13360 5900 13420
rect 5960 13360 6000 13420
rect 4460 13160 4560 13180
rect 4460 13100 4480 13160
rect 4540 13100 4560 13160
rect 1500 10780 1540 10840
rect 1600 10780 1620 10840
rect 1500 9580 1620 10780
rect 1500 9520 1540 9580
rect 1600 9520 1620 9580
rect 1879 9780 2001 11097
rect 2260 11080 2300 11140
rect 2360 11080 2380 11140
rect 2260 11060 2380 11080
rect 2920 11160 3040 11180
rect 2920 11100 2940 11160
rect 3000 11100 3040 11160
rect 1879 9720 1920 9780
rect 1980 9720 2001 9780
rect 1879 9579 2001 9720
rect 2640 9780 2740 9800
rect 2640 9720 2660 9780
rect 2720 9720 2740 9780
rect 2260 9580 2380 9600
rect 1500 8600 1620 9520
rect 1880 8620 2000 9579
rect 2260 9520 2280 9580
rect 2340 9520 2380 9580
rect 2260 8620 2380 9520
rect 2640 8620 2740 9720
rect 2920 9220 3040 11100
rect 3660 11160 3800 11180
rect 3660 11100 3700 11160
rect 3760 11100 3800 11160
rect 3280 10660 3400 10680
rect 3280 10600 3300 10660
rect 3360 10600 3400 10660
rect 3280 8620 3400 10600
rect 3660 8620 3800 11100
rect 4040 10660 4160 10680
rect 4040 10600 4080 10660
rect 4140 10600 4160 10660
rect 4040 8620 4160 10600
rect 4240 10360 4340 10380
rect 4240 10300 4260 10360
rect 4320 10300 4340 10360
rect 4240 10180 4340 10300
rect 4460 10360 4560 13100
rect 5280 12380 5340 13260
rect 5880 13120 6000 13360
rect 5880 13060 5920 13120
rect 5980 13060 6000 13120
rect 4820 10860 4940 10880
rect 4820 10800 4840 10860
rect 4900 10800 4940 10860
rect 4820 10760 4940 10800
rect 4460 10300 4480 10360
rect 4540 10300 4560 10360
rect 4460 10280 4560 10300
rect 4640 10360 4740 10380
rect 4640 10300 4660 10360
rect 4720 10300 4740 10360
rect 4640 10180 4740 10300
rect 1700 8460 1800 8560
rect 1700 8400 1720 8460
rect 1780 8400 1800 8460
rect 1700 8380 1800 8400
rect 2080 8460 2180 8560
rect 2080 8400 2100 8460
rect 2160 8400 2180 8460
rect 2080 8380 2180 8400
rect 2460 8460 2560 8560
rect 2460 8400 2480 8460
rect 2540 8400 2560 8460
rect 2460 8380 2560 8400
rect 3100 8460 3200 8560
rect 3100 8400 3120 8460
rect 3180 8400 3200 8460
rect 3100 8380 3200 8400
rect 3480 8460 3580 8560
rect 3480 8400 3500 8460
rect 3560 8400 3580 8460
rect 3480 8380 3580 8400
rect 3860 8460 3960 8560
rect 3860 8400 3880 8460
rect 3940 8400 3960 8460
rect 3860 8380 3960 8400
rect 4420 8360 4560 10120
rect 4840 9960 4940 10760
rect 5280 9500 5360 11500
rect 5880 10240 6000 13060
rect 6300 13120 6420 13140
rect 6300 13060 6320 13120
rect 6380 13060 6420 13120
rect 6300 12940 6420 13060
rect 6500 12880 6600 13580
rect 7260 13640 7360 13660
rect 7260 13580 7280 13640
rect 7340 13580 7360 13640
rect 6680 13120 6800 13140
rect 6680 13060 6700 13120
rect 6760 13060 6800 13120
rect 6680 12940 6800 13060
rect 7060 13120 7180 13140
rect 7060 13060 7080 13120
rect 7140 13060 7180 13120
rect 7060 12940 7180 13060
rect 7260 12880 7360 13580
rect 7440 13120 7560 13140
rect 7440 13060 7460 13120
rect 7520 13060 7560 13120
rect 7440 12940 7560 13060
rect 5880 10180 5920 10240
rect 5980 10180 6000 10240
rect 5880 10160 6000 10180
rect 5260 9480 5380 9500
rect 5260 9400 5280 9480
rect 5360 9400 5380 9480
rect 5260 9380 5380 9400
rect 5179 8879 5291 9154
rect 5179 8478 5185 8879
rect 5285 8478 5291 8879
rect 5179 8360 5291 8478
rect 4420 8320 5291 8360
rect 4420 8260 4460 8320
rect 4520 8260 5291 8320
rect 4420 8240 5291 8260
rect 6120 8340 6220 11800
rect 6480 10400 6620 12880
rect 6860 10400 7000 12880
rect 7240 10400 7380 12880
rect 6300 10240 6420 10340
rect 6300 10180 6320 10240
rect 6380 10180 6420 10240
rect 6300 10160 6420 10180
rect 6680 10240 6800 10340
rect 6680 10180 6700 10240
rect 6760 10180 6800 10240
rect 6680 10160 6800 10180
rect 6120 8280 6140 8340
rect 6200 8280 6220 8340
rect 6120 8240 6220 8280
rect 6880 8340 6980 10400
rect 7060 10240 7180 10340
rect 7060 10180 7080 10240
rect 7140 10180 7180 10240
rect 7060 10160 7180 10180
rect 7440 10240 7560 10340
rect 7440 10180 7460 10240
rect 7520 10180 7560 10240
rect 7440 10160 7560 10180
rect 6880 8280 6900 8340
rect 6960 8280 6980 8340
rect 6880 8240 6980 8280
rect 7640 8340 7740 11800
rect 7640 8280 7660 8340
rect 7720 8280 7740 8340
rect 7640 8240 7740 8280
rect 5179 8203 5291 8240
<< via1 >>
rect 1680 16420 1740 16480
rect 200 15800 252 15852
rect 600 15800 652 15852
rect 20 13760 80 13820
rect -360 13040 -308 13092
rect 980 15960 1032 16012
rect 2400 15960 2452 16012
rect 1340 15800 1392 15852
rect 1680 15800 1740 15860
rect 2000 15800 2052 15852
rect 780 13760 840 13820
rect 2760 15800 2812 15852
rect 3140 15800 3192 15852
rect 2580 13760 2640 13820
rect 3520 15800 3572 15852
rect 3340 13760 3400 13820
rect 2960 13580 3020 13640
rect 3720 13580 3780 13640
rect 6520 13580 6580 13640
rect 1840 13360 1900 13420
rect 2300 13360 2360 13420
rect 400 13020 452 13072
rect -560 11040 -508 11092
rect -360 11020 -300 11080
rect -180 11040 -128 11092
rect -760 10600 -700 10660
rect 1540 13100 1600 13160
rect 1920 13100 1980 13160
rect 1160 13020 1212 13072
rect 200 11040 252 11092
rect 580 11040 632 11092
rect 960 11040 1012 11092
rect 1180 11020 1240 11080
rect 1340 11040 1392 11092
rect 780 10780 840 10840
rect 0 10600 60 10660
rect -360 10380 -300 10440
rect 1180 10220 1240 10280
rect 5280 13340 5340 13400
rect 5900 13360 5960 13420
rect 4480 13100 4540 13160
rect 1540 10780 1600 10840
rect 1540 9520 1600 9580
rect 2300 11080 2360 11140
rect 2940 11100 3000 11160
rect 1920 9720 1980 9780
rect 2660 9720 2720 9780
rect 2280 9520 2340 9580
rect 3700 11100 3760 11160
rect 3300 10600 3360 10660
rect 4080 10600 4140 10660
rect 4260 10300 4320 10360
rect 5920 13060 5980 13120
rect 4840 10800 4900 10860
rect 4480 10300 4540 10360
rect 4660 10300 4720 10360
rect 1720 8400 1780 8460
rect 2100 8400 2160 8460
rect 2480 8400 2540 8460
rect 3120 8400 3180 8460
rect 3500 8400 3560 8460
rect 3880 8400 3940 8460
rect 6320 13060 6380 13120
rect 7280 13580 7340 13640
rect 6700 13060 6760 13120
rect 7080 13060 7140 13120
rect 7460 13060 7520 13120
rect 5920 10180 5980 10240
rect 5280 9400 5360 9480
rect 4460 8260 4520 8320
rect 6320 10180 6380 10240
rect 6700 10180 6760 10240
rect 6140 8280 6200 8340
rect 7080 10180 7140 10240
rect 7460 10180 7520 10240
rect 6900 8280 6960 8340
rect 7660 8280 7720 8340
<< metal2 >>
rect 1660 16480 1760 16500
rect 400 16179 460 16472
rect 1660 16420 1680 16480
rect 1740 16420 1760 16480
rect 1660 16400 1760 16420
rect 400 16119 3015 16179
rect 200 15860 252 15862
rect 400 15860 460 16119
rect 1607 16040 1667 16119
rect 960 16012 2460 16040
rect 960 15960 980 16012
rect 1032 15960 2400 16012
rect 2452 15960 2460 16012
rect 960 15940 2460 15960
rect 600 15860 652 15862
rect 1340 15860 1392 15862
rect 1680 15860 1740 15870
rect 2000 15860 2052 15862
rect 2760 15860 2812 15862
rect 2955 15860 3015 16119
rect 3140 15860 3192 15862
rect 3520 15860 3572 15862
rect 160 15852 680 15860
rect 160 15800 200 15852
rect 252 15800 600 15852
rect 652 15800 680 15852
rect 1300 15852 1680 15860
rect 1300 15800 1340 15852
rect 1392 15800 1680 15852
rect 1740 15852 2100 15860
rect 1740 15800 2000 15852
rect 2052 15800 2100 15852
rect 2720 15852 3620 15860
rect 2720 15800 2760 15852
rect 2812 15800 3140 15852
rect 3192 15800 3520 15852
rect 3572 15800 3620 15852
rect 200 15790 252 15800
rect 600 15790 652 15800
rect 1340 15790 1392 15800
rect 1680 15790 1740 15800
rect 2000 15790 2052 15800
rect 2760 15790 2812 15800
rect 3140 15790 3192 15800
rect 3520 15790 3572 15800
rect -20 13820 3420 13840
rect -20 13760 20 13820
rect 80 13760 780 13820
rect 840 13760 2580 13820
rect 2640 13760 3340 13820
rect 3400 13760 3420 13820
rect -20 13740 3420 13760
rect 4780 13660 4880 16500
rect 2920 13640 8030 13660
rect 2920 13580 2960 13640
rect 3020 13580 3720 13640
rect 3780 13580 6520 13640
rect 6580 13580 7280 13640
rect 7340 13580 7960 13640
rect 8020 13580 8030 13640
rect 2920 13560 8030 13580
rect 1800 13420 6000 13440
rect 1800 13360 1840 13420
rect 1900 13360 2300 13420
rect 2360 13400 5900 13420
rect 2360 13360 5280 13400
rect 1800 13340 5280 13360
rect 5340 13360 5900 13400
rect 5960 13360 6000 13420
rect 5340 13340 6000 13360
rect 1800 13320 6000 13340
rect 1500 13160 4560 13180
rect -400 13092 1240 13120
rect -400 13040 -360 13092
rect -308 13072 1240 13092
rect 1500 13100 1540 13160
rect 1600 13100 1920 13160
rect 1980 13100 4480 13160
rect 4540 13100 4560 13160
rect 1500 13080 4560 13100
rect 5880 13120 7560 13140
rect -308 13040 400 13072
rect -400 13020 400 13040
rect 452 13020 1160 13072
rect 1212 13020 1240 13072
rect 5880 13060 5920 13120
rect 5980 13060 6320 13120
rect 6380 13060 6700 13120
rect 6760 13060 7080 13120
rect 7140 13060 7460 13120
rect 7520 13060 7560 13120
rect 5880 13040 7560 13060
rect -400 12980 1240 13020
rect 2260 11160 3800 11180
rect 2260 11140 2940 11160
rect -560 11100 -508 11102
rect -180 11100 -128 11102
rect 200 11100 252 11102
rect 580 11100 632 11102
rect 960 11100 1012 11102
rect 1340 11100 1392 11102
rect -580 11092 280 11100
rect -580 11040 -560 11092
rect -508 11080 -180 11092
rect -508 11040 -360 11080
rect -580 11020 -360 11040
rect -300 11040 -180 11080
rect -128 11040 200 11092
rect 252 11040 280 11092
rect -300 11020 280 11040
rect 560 11092 1420 11100
rect 560 11040 580 11092
rect 632 11040 960 11092
rect 1012 11080 1340 11092
rect 1012 11040 1180 11080
rect 560 11020 1180 11040
rect 1240 11040 1340 11080
rect 1392 11040 1420 11092
rect 2260 11080 2300 11140
rect 2360 11100 2940 11140
rect 3000 11100 3700 11160
rect 3760 11100 3800 11160
rect 2360 11080 3800 11100
rect 2260 11060 3800 11080
rect 1240 11020 1420 11040
rect -360 11010 -300 11020
rect 1180 11010 1240 11020
rect 740 10860 4940 10880
rect 740 10840 4840 10860
rect 740 10780 780 10840
rect 840 10780 1540 10840
rect 1600 10800 4840 10840
rect 4900 10800 4940 10860
rect 1600 10780 4940 10800
rect 740 10760 4940 10780
rect -800 10660 4160 10680
rect -800 10600 -760 10660
rect -700 10600 0 10660
rect 60 10600 3300 10660
rect 3360 10600 4080 10660
rect 4140 10600 4160 10660
rect -800 10580 4160 10600
rect -1320 10440 -280 10460
rect -1320 10380 -360 10440
rect -300 10380 -280 10440
rect -1320 10360 -280 10380
rect 4240 10360 4740 10380
rect 4240 10300 4260 10360
rect 4320 10300 4480 10360
rect 4540 10300 4660 10360
rect 4720 10300 4740 10360
rect -1320 10280 1280 10300
rect 4240 10280 4740 10300
rect -1320 10220 1180 10280
rect 1240 10220 1280 10280
rect -1320 10200 1280 10220
rect 5880 10240 7560 10260
rect 5880 10180 5920 10240
rect 5980 10180 6320 10240
rect 6380 10180 6700 10240
rect 6760 10180 7080 10240
rect 7140 10180 7460 10240
rect 7520 10180 7560 10240
rect 5880 10160 7560 10180
rect 1880 9780 2740 9800
rect 1880 9720 1920 9780
rect 1980 9720 2660 9780
rect 2720 9720 2740 9780
rect 1880 9700 2740 9720
rect 1500 9580 2380 9600
rect 1500 9520 1540 9580
rect 1600 9520 2280 9580
rect 2340 9520 2380 9580
rect 1500 9500 2380 9520
rect 5260 9480 5380 9500
rect 5260 9400 5280 9480
rect 5360 9400 5380 9480
rect 5260 9380 5380 9400
rect -1320 8460 3960 8480
rect -1320 8400 1720 8460
rect 1780 8400 2100 8460
rect 2160 8400 2480 8460
rect 2540 8400 3120 8460
rect 3180 8400 3500 8460
rect 3560 8400 3880 8460
rect 3940 8400 3960 8460
rect -1320 8380 3960 8400
rect 4420 8340 7740 8360
rect 4420 8320 6140 8340
rect 4420 8260 4460 8320
rect 4520 8280 6140 8320
rect 6200 8280 6900 8340
rect 6960 8280 7660 8340
rect 7720 8280 7740 8340
rect 4520 8260 7740 8280
rect 4420 8240 7740 8260
rect 4820 7800 4920 8240
<< via2 >>
rect 7960 13580 8020 13640
rect 5280 9400 5360 9480
<< metal3 >>
rect 7940 13640 8060 13660
rect 7940 13580 7960 13640
rect 8020 13580 8060 13640
rect 7940 13080 8060 13580
rect 7940 13000 7960 13080
rect 8040 13000 8060 13080
rect 7940 12980 8060 13000
rect 5260 9480 5380 9500
rect 5260 9400 5280 9480
rect 5360 9400 5380 9480
rect 5260 9380 5380 9400
<< via3 >>
rect 7960 13000 8040 13080
rect 5280 9400 5360 9480
<< metal4 >>
rect 8080 13160 8520 13260
rect 8080 13100 8160 13160
rect 7940 13080 8160 13100
rect 7940 13000 7960 13080
rect 8040 13000 8160 13080
rect 7940 12980 8160 13000
rect 8080 12920 8160 12980
rect 8400 12920 8520 13160
rect 8080 12820 8520 12920
rect 8160 9560 8560 9660
rect 8160 9500 8240 9560
rect 5260 9480 8240 9500
rect 5260 9400 5280 9480
rect 5360 9400 8240 9480
rect 5260 9380 8240 9400
rect 8160 9320 8240 9380
rect 8480 9320 8560 9560
rect 8160 9220 8560 9320
<< via4 >>
rect 8160 12920 8400 13160
rect 8240 9320 8480 9560
<< metal5 >>
rect 8080 13160 9060 13260
rect 8080 12920 8160 13160
rect 8400 12920 9060 13160
rect 8080 12820 9060 12920
rect 10040 9660 10360 10320
rect 8160 9560 10360 9660
rect 8160 9320 8240 9560
rect 8480 9320 10360 9560
rect 8160 9220 10360 9320
use sky130_fd_pr__nfet_01v8_7JHNGK  sky130_fd_pr__nfet_01v8_7JHNGK_0
timestamp 1733707933
transform 1 0 4698 0 1 9377
box -158 -857 158 857
use sky130_fd_pr__nfet_01v8_7JHNGK  sky130_fd_pr__nfet_01v8_7JHNGK_1
timestamp 1733707933
transform 1 0 4298 0 1 9377
box -158 -857 158 857
use sky130_fd_pr__nfet_01v8_Q7LUJ6  sky130_fd_pr__nfet_01v8_Q7LUJ6_0
timestamp 1733700048
transform 1 0 7498 0 1 10957
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7LUJ6  sky130_fd_pr__nfet_01v8_Q7LUJ6_1
timestamp 1733700048
transform 1 0 6358 0 1 10957
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7LUJ6  sky130_fd_pr__nfet_01v8_Q7LUJ6_2
timestamp 1733700048
transform 1 0 6738 0 1 10957
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7LUJ6  sky130_fd_pr__nfet_01v8_Q7LUJ6_3
timestamp 1733700048
transform 1 0 7118 0 1 10957
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7ZM59  sky130_fd_pr__nfet_01v8_Q7ZM59_0
timestamp 1733700048
transform 1 0 7118 0 1 12317
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7ZM59  sky130_fd_pr__nfet_01v8_Q7ZM59_1
timestamp 1733700048
transform 1 0 7498 0 1 12317
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7ZM59  sky130_fd_pr__nfet_01v8_Q7ZM59_2
timestamp 1733700048
transform 1 0 6358 0 1 12317
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_Q7ZM59  sky130_fd_pr__nfet_01v8_Q7ZM59_3
timestamp 1733700048
transform 1 0 6738 0 1 12317
box -158 -657 158 657
use sky130_fd_pr__nfet_01v8_QP3KE5  sky130_fd_pr__nfet_01v8_QP3KE5_0
timestamp 1733700048
transform -1 0 2518 0 -1 8977
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_QP3KE5  sky130_fd_pr__nfet_01v8_QP3KE5_1
timestamp 1733700048
transform -1 0 1758 0 -1 8977
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_QP3KE5  sky130_fd_pr__nfet_01v8_QP3KE5_2
timestamp 1733700048
transform -1 0 2138 0 -1 8977
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_QP3KE5  sky130_fd_pr__nfet_01v8_QP3KE5_3
timestamp 1733700048
transform -1 0 3538 0 -1 8977
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_QP3KE5  sky130_fd_pr__nfet_01v8_QP3KE5_4
timestamp 1733700048
transform -1 0 3158 0 -1 8977
box -158 -457 158 457
use sky130_fd_pr__nfet_01v8_QP3KE5  sky130_fd_pr__nfet_01v8_QP3KE5_5
timestamp 1733700048
transform -1 0 3918 0 -1 8977
box -158 -457 158 457
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_0
timestamp 1733715709
transform 1 0 234 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_1
timestamp 1733715709
transform 1 0 614 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_2
timestamp 1733715709
transform 1 0 994 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_3
timestamp 1733715709
transform 1 0 1374 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_4
timestamp 1733715709
transform 1 0 2034 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_5
timestamp 1733715709
transform 1 0 2414 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_6
timestamp 1733715709
transform 1 0 2794 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_7
timestamp 1733715709
transform 1 0 3174 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_EXDZWJ  sky130_fd_pr__pfet_01v8_lvt_EXDZWJ_8
timestamp 1733715709
transform 1 0 3554 0 1 14898
box -194 -998 194 964
use sky130_fd_pr__pfet_01v8_lvt_NBBSEP  sky130_fd_pr__pfet_01v8_lvt_NBBSEP_0
timestamp 1733715709
transform -1 0 994 0 -1 12044
box -194 -898 194 864
use sky130_fd_pr__pfet_01v8_lvt_NBBSEP  sky130_fd_pr__pfet_01v8_lvt_NBBSEP_1
timestamp 1733715709
transform -1 0 -526 0 -1 12044
box -194 -898 194 864
use sky130_fd_pr__pfet_01v8_lvt_NBBSEP  sky130_fd_pr__pfet_01v8_lvt_NBBSEP_2
timestamp 1733715709
transform -1 0 -146 0 -1 12044
box -194 -898 194 864
use sky130_fd_pr__pfet_01v8_lvt_NBBSEP  sky130_fd_pr__pfet_01v8_lvt_NBBSEP_3
timestamp 1733715709
transform -1 0 234 0 -1 12044
box -194 -898 194 864
use sky130_fd_pr__pfet_01v8_lvt_NBBSEP  sky130_fd_pr__pfet_01v8_lvt_NBBSEP_4
timestamp 1733715709
transform -1 0 1374 0 -1 12044
box -194 -898 194 864
use sky130_fd_pr__pfet_01v8_lvt_NXDZEP  sky130_fd_pr__pfet_01v8_lvt_NXDZEP_0
timestamp 1733715975
transform -1 0 614 0 -1 12044
box -194 -898 194 864
use sky130_fd_pr__res_xhigh_po_0p35_QT585A  sky130_fd_pr__res_xhigh_po_0p35_QT585A_0
timestamp 1733710384
transform 1 0 5315 0 1 11982
box -35 -542 35 542
use sky130_fd_pr__cap_mim_m3_2_KAF84V  XC2
timestamp 1733700048
transform -1 0 9931 0 -1 13860
box -1049 -3600 1071 3600
<< labels >>
rlabel metal2 400 16412 460 16472 1 Vb1
port 1 n
rlabel metal2 -1300 10220 -1240 10280 1 Vinm
port 2 n
rlabel metal2 -1300 10380 -1240 10440 1 Vinp
port 3 n
rlabel metal2 1680 16420 1740 16480 1 Vb2
port 4 n
rlabel metal2 -1300 8400 -1240 8460 1 Vb3
port 5 n
rlabel metal2 4800 16420 4860 16480 1 Vout
port 6 n
rlabel metal1 -1220 15540 -1160 15600 1 VDD
port 7 n
rlabel metal2 4840 7820 4900 7880 1 VSS
port 8 n
<< properties >>
string FIXED_BBOX -9872 928 1812 7312
<< end >>
