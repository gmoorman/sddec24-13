magic
tech sky130B
magscale 1 2
timestamp 1733710384
<< xpolycontact >>
rect -35 110 35 542
rect -35 -542 35 -110
<< xpolyres >>
rect -35 -110 35 110
<< viali >>
rect -19 127 19 524
rect -19 -524 19 -127
<< metal1 >>
rect -25 524 25 536
rect -25 127 -19 524
rect 19 127 25 524
rect -25 115 25 127
rect -25 -127 25 -115
rect -25 -524 -19 -127
rect 19 -524 25 -127
rect -25 -536 25 -524
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.1 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 7.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
