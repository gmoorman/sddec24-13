magic
tech sky130B
magscale 1 2
timestamp 1733695688
<< pwell >>
rect -201 -1362 201 1362
<< psubdiff >>
rect -165 1292 -69 1326
rect 69 1292 165 1326
rect -165 1230 -131 1292
rect 131 1230 165 1292
rect -165 -1292 -131 -1230
rect 131 -1292 165 -1230
rect -165 -1326 -69 -1292
rect 69 -1326 165 -1292
<< psubdiffcont >>
rect -69 1292 69 1326
rect -165 -1230 -131 1230
rect 131 -1230 165 1230
rect -69 -1326 69 -1292
<< xpolycontact >>
rect -35 764 35 1196
rect -35 52 35 484
rect -35 -484 35 -52
rect -35 -1196 35 -764
<< xpolyres >>
rect -35 484 35 764
rect -35 -764 35 -484
<< locali >>
rect -165 1292 -69 1326
rect 69 1292 165 1326
rect -165 1230 -131 1292
rect 131 1230 165 1292
rect -165 -1292 -131 -1230
rect 131 -1292 165 -1230
rect -165 -1326 -69 -1292
rect 69 -1326 165 -1292
<< viali >>
rect -19 781 19 1178
rect -19 70 19 467
rect -19 -467 19 -70
rect -19 -1178 19 -781
<< metal1 >>
rect -25 1178 25 1190
rect -25 781 -19 1178
rect 19 781 25 1178
rect -25 769 25 781
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect -25 -781 25 -769
rect -25 -1178 -19 -781
rect 19 -1178 25 -781
rect -25 -1190 25 -1178
<< properties >>
string FIXED_BBOX -148 -1309 148 1309
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.562 m 2 nx 1 wmin 0.350 lmin 0.50 class resistor rho 2000 val 10.001k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
