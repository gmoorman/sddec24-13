magic
tech sky130B
magscale 1 2
timestamp 1733695688
<< pwell >>
rect -201 -738 201 738
<< psubdiff >>
rect -165 668 -69 702
rect 69 668 165 702
rect -165 606 -131 668
rect 131 606 165 668
rect -165 -668 -131 -606
rect 131 -668 165 -606
rect -165 -702 -69 -668
rect 69 -702 165 -668
<< psubdiffcont >>
rect -69 668 69 702
rect -165 -606 -131 606
rect 131 -606 165 606
rect -69 -702 69 -668
<< xpolycontact >>
rect -35 140 35 572
rect -35 -572 35 -140
<< xpolyres >>
rect -35 -140 35 140
<< locali >>
rect -165 668 -69 702
rect 69 668 165 702
rect -165 606 -131 668
rect 131 606 165 668
rect -165 -668 -131 -606
rect 131 -668 165 -606
rect -165 -702 -69 -668
rect 69 -702 165 -668
<< viali >>
rect -19 157 19 554
rect -19 -554 19 -157
<< metal1 >>
rect -25 554 25 566
rect -25 157 -19 554
rect 19 157 25 554
rect -25 145 25 157
rect -25 -157 25 -145
rect -25 -554 -19 -157
rect 19 -554 25 -157
rect -25 -566 25 -554
<< properties >>
string FIXED_BBOX -148 -685 148 685
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.562 m 1 nx 1 wmin 0.350 lmin 0.50 class resistor rho 2000 val 10.001k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
