magic
tech sky130B
magscale 1 2
timestamp 1732510450
<< pwell >>
rect -574 -8600 3812 -1900
<< mvpsubdiff >>
rect -508 -1978 3746 -1966
rect -508 -2078 -334 -1978
rect 3572 -2078 3746 -1978
rect -508 -2090 3746 -2078
rect -508 -2140 -384 -2090
rect -508 -8360 -496 -2140
rect -396 -8360 -384 -2140
rect -508 -8410 -384 -8360
rect 3622 -2140 3746 -2090
rect 3622 -8360 3634 -2140
rect 3734 -8360 3746 -2140
rect 3622 -8410 3746 -8360
rect -508 -8422 3746 -8410
rect -508 -8522 -334 -8422
rect 3572 -8522 3746 -8422
rect -508 -8534 3746 -8522
<< mvpsubdiffcont >>
rect -334 -2078 3572 -1978
rect -496 -8360 -396 -2140
rect 3634 -8360 3734 -2140
rect -334 -8522 3572 -8422
<< locali >>
rect -496 -2140 -396 -1978
rect -496 -8522 -396 -8360
rect 3634 -2140 3734 -1978
rect 3634 -8522 3734 -8360
<< viali >>
rect -396 -2078 -334 -1978
rect -334 -2078 3572 -1978
rect 3572 -2078 3634 -1978
rect -496 -8105 -396 -2395
rect 3634 -8105 3734 -2395
rect -396 -8522 -334 -8422
rect -334 -8522 3572 -8422
rect 3572 -8522 3634 -8422
<< metal1 >>
rect -502 -1978 3740 -1972
rect -502 -2078 -396 -1978
rect 3634 -2078 3740 -1978
rect -502 -2084 3740 -2078
rect -502 -2395 -390 -2084
rect -502 -8105 -496 -2395
rect -396 -8105 -390 -2395
rect -502 -8416 -390 -8105
rect 3628 -2395 3740 -2084
rect 3628 -8105 3634 -2395
rect 3734 -8105 3740 -2395
rect 210 -8416 220 -8116
rect 3018 -8416 3028 -8116
rect 3628 -8416 3740 -8105
rect -502 -8422 3740 -8416
rect -502 -8522 -396 -8422
rect 3634 -8522 3740 -8422
rect -502 -8528 3740 -8522
<< via1 >>
rect -390 -8416 210 -8116
rect 3028 -8416 3628 -8116
<< metal2 >>
rect -390 -8116 210 -8106
rect -390 -8426 210 -8416
rect 3028 -8116 3628 -8106
rect 3028 -8426 3628 -8416
<< via2 >>
rect -390 -8416 210 -8116
rect 3028 -8416 3628 -8116
<< metal3 >>
rect -400 -8116 220 -8111
rect -400 -8416 -390 -8116
rect 210 -8416 220 -8116
rect -400 -8421 220 -8416
rect 3018 -8116 3638 -8111
rect 3018 -8416 3028 -8116
rect 3628 -8416 3638 -8116
rect 3018 -8421 3638 -8416
<< via3 >>
rect -390 -8416 210 -8116
rect 3028 -8416 3628 -8116
<< metal4 >>
rect -391 -8116 211 -8115
rect -391 -8416 -390 -8116
rect 210 -8416 211 -8116
rect -391 -8417 211 -8416
rect 3027 -8116 3629 -8115
rect 3027 -8416 3028 -8116
rect 3628 -8416 3629 -8116
rect 3027 -8417 3629 -8416
<< properties >>
string FIXED_BBOX -446 -8472 3684 -2028
<< end >>
