magic
tech sky130B
magscale 1 2
timestamp 1733645871
<< nwell >>
rect -574 -1788 3812 1200
<< pwell >>
rect -574 -8600 3812 -1900
<< mvpsubdiff >>
rect -508 -1978 3746 -1966
rect -508 -2078 -334 -1978
rect 3572 -2078 3746 -1978
rect -508 -2090 3746 -2078
rect -508 -2140 -384 -2090
rect -508 -8360 -496 -2140
rect -396 -8360 -384 -2140
rect -508 -8410 -384 -8360
rect 3622 -2140 3746 -2090
rect 3622 -8360 3634 -2140
rect 3734 -8360 3746 -2140
rect 3622 -8410 3746 -8360
rect -508 -8422 3746 -8410
rect -508 -8522 -334 -8422
rect 3572 -8522 3746 -8422
rect -508 -8534 3746 -8522
<< mvnsubdiff >>
rect -508 1122 3746 1134
rect -508 1022 -334 1122
rect 3572 1022 3746 1122
rect -508 1010 3746 1022
rect -508 960 -384 1010
rect -508 -1548 -496 960
rect -396 -1548 -384 960
rect -508 -1598 -384 -1548
rect 3622 960 3746 1010
rect 3622 -1548 3634 960
rect 3734 -1548 3746 960
rect 3622 -1598 3746 -1548
rect -508 -1610 3746 -1598
rect -508 -1710 -334 -1610
rect 3572 -1710 3746 -1610
rect -508 -1722 3746 -1710
<< mvpsubdiffcont >>
rect -334 -2078 3572 -1978
rect -496 -8360 -396 -2140
rect 3634 -8360 3734 -2140
rect -334 -8522 3572 -8422
<< mvnsubdiffcont >>
rect -334 1022 3572 1122
rect -496 -1548 -396 960
rect 3634 -1548 3734 960
rect -334 -1710 3572 -1610
<< locali >>
rect -496 960 -396 1122
rect -496 -1710 -396 -1548
rect 3634 960 3734 1122
rect 3634 -1710 3734 -1548
rect -496 -2140 -396 -1978
rect -496 -8522 -396 -8360
rect 3634 -2140 3734 -1978
rect 3634 -8522 3734 -8360
<< viali >>
rect -396 1022 -334 1122
rect -334 1022 3572 1122
rect 3572 1022 3634 1122
rect -496 -1478 -396 890
rect 3634 -1478 3734 890
rect -396 -1710 -334 -1610
rect -334 -1710 3572 -1610
rect 3572 -1710 3634 -1610
rect -396 -2078 -334 -1978
rect -334 -2078 3572 -1978
rect 3572 -2078 3634 -1978
rect -496 -8105 -396 -2395
rect 3634 -8105 3734 -2395
rect -396 -8522 -334 -8422
rect -334 -8522 3572 -8422
rect 3572 -8522 3634 -8422
<< metal1 >>
rect -502 1122 3740 1128
rect -502 1022 -396 1122
rect 3634 1022 3740 1122
rect -502 1016 3740 1022
rect -502 890 -390 1016
rect -502 -1478 -496 890
rect -396 -1478 -390 890
rect 210 716 220 1016
rect 3018 716 3028 1016
rect 3628 890 3740 1016
rect -110 492 -58 716
rect -110 -684 -58 440
rect 170 492 222 502
rect -26 398 26 408
rect -26 336 26 346
rect -18 246 18 336
rect -18 -308 18 -246
rect 60 -330 112 -30
rect -18 -470 18 -408
rect -18 -1052 18 -962
rect -26 -1062 26 -1052
rect -26 -1124 26 -1114
rect 60 -1300 112 -382
rect 170 -684 222 440
rect 450 492 502 502
rect 254 398 306 408
rect 254 336 306 346
rect 262 246 298 336
rect 262 -308 298 -246
rect 340 -330 392 -30
rect 262 -470 298 -408
rect 340 -682 392 -382
rect 450 -684 502 440
rect 730 492 782 498
rect 534 398 586 408
rect 534 336 586 346
rect 542 246 578 336
rect 542 -308 578 -246
rect 620 -330 672 -30
rect 542 -470 578 -408
rect 620 -682 672 -382
rect 730 -684 782 440
rect 1010 492 1062 502
rect 814 398 866 408
rect 814 336 866 346
rect 822 246 858 336
rect 822 -308 858 -246
rect 900 -330 952 -30
rect 822 -470 858 -408
rect 900 -682 952 -382
rect 1010 -684 1062 440
rect 1290 492 1342 502
rect 1094 398 1146 408
rect 1094 336 1146 346
rect 1102 246 1138 336
rect 1102 -308 1138 -246
rect 1180 -330 1232 -30
rect 1102 -470 1138 -408
rect 1180 -682 1232 -382
rect 1290 -684 1342 440
rect 1570 492 1622 502
rect 1374 398 1426 408
rect 1374 336 1426 346
rect 1382 246 1418 336
rect 1382 -308 1418 -246
rect 1460 -330 1512 -30
rect 1382 -470 1418 -408
rect 1460 -682 1512 -382
rect 1570 -684 1622 440
rect 1850 492 1902 502
rect 1654 398 1706 408
rect 1654 336 1706 346
rect 1662 246 1698 336
rect 1662 -308 1698 -246
rect 1740 -330 1792 -30
rect 1662 -470 1698 -408
rect 1740 -682 1792 -382
rect 1850 -684 1902 440
rect 2130 492 2182 502
rect 1934 398 1986 408
rect 1934 336 1986 346
rect 1942 246 1978 336
rect 1942 -308 1978 -246
rect 2020 -330 2072 -30
rect 1942 -470 1978 -408
rect 2020 -682 2072 -382
rect 2130 -684 2182 440
rect 2410 492 2462 502
rect 2214 398 2266 408
rect 2214 336 2266 346
rect 2222 246 2258 336
rect 2222 -308 2258 -246
rect 2300 -330 2352 -30
rect 2222 -470 2258 -408
rect 2300 -682 2352 -382
rect 2410 -684 2462 440
rect 2690 492 2742 502
rect 2494 398 2546 408
rect 2494 336 2546 346
rect 2502 246 2538 336
rect 2502 -308 2538 -246
rect 2580 -330 2632 -30
rect 2502 -470 2538 -408
rect 2580 -682 2632 -382
rect 2690 -684 2742 440
rect 2970 492 3022 502
rect 2774 398 2826 408
rect 2774 336 2826 346
rect 2782 246 2818 336
rect 2782 -308 2818 -246
rect 2860 -330 2912 -30
rect 2782 -470 2818 -408
rect 2860 -682 2912 -382
rect 2970 -684 3022 440
rect 3228 282 3238 290
rect 3062 246 3238 282
rect 3228 238 3238 246
rect 3290 238 3520 290
rect 3572 238 3582 290
rect 3062 -308 3098 -246
rect 3140 -330 3192 -30
rect 3062 -470 3098 -408
rect 262 -1052 298 -962
rect 542 -1052 578 -962
rect 822 -1052 858 -962
rect 1102 -1052 1138 -962
rect 254 -1062 306 -1052
rect 254 -1124 306 -1114
rect 534 -1062 586 -1052
rect 534 -1124 586 -1114
rect 814 -1062 866 -1052
rect 814 -1124 866 -1114
rect 1094 -1062 1146 -1052
rect 1094 -1124 1146 -1114
rect 1382 -1168 1418 -962
rect 1662 -1168 1698 -962
rect 1942 -1052 1978 -962
rect 2222 -1052 2258 -962
rect 2502 -1052 2538 -962
rect 2782 -1052 2818 -962
rect 3062 -1052 3098 -962
rect 1934 -1062 1986 -1052
rect 1934 -1124 1986 -1114
rect 2214 -1062 2266 -1052
rect 2214 -1124 2266 -1114
rect 2494 -1062 2546 -1052
rect 2494 -1124 2546 -1114
rect 2774 -1062 2826 -1052
rect 2774 -1124 2826 -1114
rect 3054 -1062 3106 -1052
rect 3054 -1124 3106 -1114
rect 1374 -1178 1426 -1168
rect 1374 -1240 1426 -1230
rect 1654 -1178 1706 -1168
rect 1654 -1240 1706 -1230
rect -502 -1604 -390 -1478
rect 66 -1472 102 -1300
rect 404 -1472 414 -1462
rect 66 -1508 414 -1472
rect 404 -1514 414 -1508
rect 466 -1472 476 -1462
rect 1662 -1472 1698 -1240
rect 3140 -1372 3192 -382
rect 2468 -1424 2478 -1372
rect 2530 -1424 3192 -1372
rect 466 -1508 1698 -1472
rect 3628 -1478 3634 890
rect 3734 -1478 3740 890
rect 466 -1514 476 -1508
rect 3628 -1604 3740 -1478
rect -502 -1610 3740 -1604
rect -502 -1710 -396 -1610
rect 3634 -1710 3740 -1610
rect -502 -1716 3740 -1710
rect -502 -1978 3740 -1972
rect -502 -2078 -396 -1978
rect 3634 -2078 3740 -1978
rect -502 -2084 3740 -2078
rect -502 -2395 -390 -2084
rect 900 -2142 952 -2132
rect 900 -2204 952 -2194
rect 2774 -2134 2826 -2124
rect 2774 -2196 2826 -2186
rect 330 -2222 382 -2212
rect 330 -2284 382 -2274
rect 610 -2222 662 -2212
rect 610 -2284 662 -2274
rect 178 -2322 230 -2312
rect 178 -2384 230 -2374
rect -502 -8105 -496 -2395
rect -396 -2742 -390 -2395
rect 186 -2670 222 -2384
rect 254 -2422 306 -2412
rect 254 -2484 306 -2474
rect 262 -2538 298 -2484
rect 338 -2670 374 -2284
rect 458 -2322 510 -2312
rect 458 -2384 510 -2374
rect 466 -2670 502 -2384
rect 534 -2422 586 -2412
rect 534 -2484 586 -2474
rect 542 -2538 578 -2484
rect 618 -2670 654 -2284
rect 814 -2422 866 -2412
rect 814 -2484 866 -2474
rect 822 -2538 858 -2484
rect -396 -2778 50 -2742
rect -396 -2984 -390 -2778
rect 900 -2950 936 -2204
rect 1450 -2222 1502 -2212
rect 1450 -2284 1502 -2274
rect 1730 -2222 1782 -2212
rect 1730 -2284 1782 -2274
rect 2570 -2222 2622 -2212
rect 2570 -2284 2622 -2274
rect 1298 -2322 1350 -2312
rect 1298 -2384 1350 -2374
rect 1094 -2422 1146 -2412
rect 1094 -2484 1146 -2474
rect 1102 -2538 1138 -2484
rect 1306 -2670 1342 -2384
rect 1374 -2422 1426 -2412
rect 1374 -2484 1426 -2474
rect 1382 -2538 1418 -2484
rect 1458 -2670 1494 -2284
rect 1578 -2322 1630 -2312
rect 1578 -2384 1630 -2374
rect 1586 -2670 1622 -2384
rect 1654 -2422 1706 -2412
rect 1654 -2484 1706 -2474
rect 1662 -2538 1698 -2484
rect 1738 -2670 1774 -2284
rect 2418 -2322 2470 -2312
rect 2418 -2384 2470 -2374
rect 1934 -2422 1986 -2412
rect 1934 -2484 1986 -2474
rect 2214 -2422 2266 -2412
rect 2214 -2484 2266 -2474
rect 1942 -2538 1978 -2484
rect 2222 -2538 2258 -2484
rect 2426 -2670 2462 -2384
rect 2494 -2422 2546 -2412
rect 2494 -2484 2546 -2474
rect 2502 -2538 2538 -2484
rect 2578 -2670 2614 -2284
rect 2698 -2322 2750 -2312
rect 2698 -2384 2750 -2374
rect 2706 -2670 2742 -2384
rect 2782 -2412 2818 -2196
rect 2850 -2222 2902 -2212
rect 2850 -2284 2902 -2274
rect 2774 -2422 2826 -2412
rect 2774 -2484 2826 -2474
rect 2782 -2538 2818 -2484
rect 2858 -2670 2894 -2284
rect 3628 -2395 3740 -2084
rect 3628 -2726 3634 -2395
rect 3044 -2762 3634 -2726
rect -396 -3020 18 -2984
rect -396 -3356 -390 -3020
rect 262 -3108 298 -3048
rect 542 -3108 578 -3048
rect 746 -3132 782 -2950
rect 822 -3108 858 -3048
rect 898 -3054 936 -2950
rect 178 -3146 230 -3136
rect 178 -3208 230 -3198
rect 458 -3146 510 -3136
rect 458 -3208 510 -3198
rect 738 -3142 790 -3132
rect 738 -3204 790 -3194
rect -396 -3392 19 -3356
rect -396 -3614 -390 -3392
rect 186 -3488 222 -3208
rect 330 -3246 382 -3236
rect 330 -3308 382 -3298
rect 262 -3392 298 -3332
rect 338 -3490 374 -3308
rect 466 -3490 502 -3208
rect 898 -3236 934 -3054
rect 1026 -3132 1062 -2950
rect 1102 -3108 1138 -3048
rect 1018 -3142 1070 -3132
rect 1018 -3204 1070 -3194
rect 1178 -3236 1214 -2950
rect 1382 -3108 1418 -3048
rect 1662 -3108 1698 -3048
rect 1866 -3132 1902 -2950
rect 1942 -3108 1978 -3048
rect 1298 -3146 1350 -3136
rect 1298 -3208 1350 -3198
rect 1578 -3146 1630 -3136
rect 1578 -3208 1630 -3198
rect 1858 -3142 1910 -3132
rect 1858 -3204 1910 -3194
rect 610 -3246 662 -3236
rect 610 -3308 662 -3298
rect 890 -3246 942 -3236
rect 890 -3308 942 -3298
rect 1170 -3246 1222 -3236
rect 1170 -3308 1222 -3298
rect 542 -3392 578 -3332
rect 618 -3490 654 -3308
rect 822 -3392 858 -3332
rect 1102 -3392 1138 -3332
rect 1306 -3490 1342 -3208
rect 1450 -3246 1502 -3236
rect 1450 -3308 1502 -3298
rect 1382 -3392 1418 -3332
rect 1458 -3490 1494 -3308
rect -396 -3652 50 -3614
rect -396 -4840 -390 -3652
rect 262 -3956 298 -3902
rect 542 -3956 578 -3902
rect 254 -3966 306 -3956
rect 254 -4028 306 -4018
rect 534 -3966 586 -3956
rect 534 -4028 586 -4018
rect 746 -4156 782 -3770
rect 822 -3956 858 -3902
rect 814 -3966 866 -3956
rect 814 -4028 866 -4018
rect 898 -4056 934 -3770
rect 890 -4066 942 -4056
rect 890 -4128 942 -4118
rect 1026 -4156 1062 -3770
rect 1102 -3956 1138 -3902
rect 1094 -3966 1146 -3956
rect 1094 -4028 1146 -4018
rect 1178 -4056 1214 -3770
rect 1382 -3956 1418 -3902
rect 1374 -3966 1426 -3956
rect 1374 -4028 1426 -4018
rect 1170 -4066 1222 -4056
rect 1170 -4128 1222 -4118
rect 738 -4166 790 -4156
rect 738 -4228 790 -4218
rect 1018 -4166 1070 -4156
rect 1018 -4228 1070 -4218
rect 1178 -4328 1212 -4128
rect 1178 -4358 1418 -4328
rect 1382 -4636 1418 -4358
rect 1586 -4390 1622 -3208
rect 2018 -3236 2054 -2950
rect 2146 -3132 2182 -2950
rect 2222 -3108 2258 -3048
rect 2138 -3142 2190 -3132
rect 2138 -3204 2190 -3194
rect 2298 -3236 2334 -2950
rect 3628 -2984 3634 -2762
rect 3062 -3020 3634 -2984
rect 2502 -3108 2538 -3048
rect 2782 -3108 2818 -3048
rect 2418 -3146 2470 -3136
rect 2418 -3208 2470 -3198
rect 2698 -3146 2750 -3136
rect 2698 -3208 2750 -3198
rect 1730 -3246 1782 -3236
rect 1730 -3308 1782 -3298
rect 2010 -3246 2062 -3236
rect 2010 -3308 2062 -3298
rect 2290 -3246 2342 -3236
rect 2290 -3308 2342 -3298
rect 1662 -3392 1698 -3332
rect 1738 -3490 1774 -3308
rect 1942 -3392 1978 -3332
rect 2222 -3392 2258 -3332
rect 2426 -3490 2462 -3208
rect 2570 -3246 2622 -3236
rect 2570 -3308 2622 -3298
rect 2502 -3392 2538 -3332
rect 2578 -3490 2614 -3308
rect 2706 -3490 2742 -3208
rect 2850 -3246 2902 -3236
rect 2850 -3308 2902 -3298
rect 2782 -3392 2818 -3332
rect 2858 -3490 2894 -3308
rect 3628 -3356 3634 -3020
rect 3060 -3392 3634 -3356
rect 1662 -3956 1698 -3902
rect 1654 -3966 1706 -3956
rect 1654 -4028 1706 -4018
rect 1740 -4246 1774 -3490
rect 3628 -3616 3634 -3392
rect 3028 -3652 3634 -3616
rect 1866 -4156 1902 -3770
rect 1942 -3956 1978 -3902
rect 1934 -3966 1986 -3956
rect 1934 -4028 1986 -4018
rect 2018 -4056 2054 -3770
rect 2010 -4066 2062 -4056
rect 2010 -4128 2062 -4118
rect 2146 -4156 2182 -3770
rect 2222 -3956 2258 -3902
rect 2214 -3966 2266 -3956
rect 2214 -4028 2266 -4018
rect 2298 -4056 2334 -3770
rect 2502 -3956 2538 -3902
rect 2782 -3956 2818 -3902
rect 2494 -3966 2546 -3956
rect 2494 -4028 2546 -4018
rect 2774 -3966 2826 -3956
rect 2774 -4028 2826 -4018
rect 2290 -4066 2342 -4056
rect 2290 -4128 2342 -4118
rect 1858 -4166 1910 -4156
rect 1858 -4228 1910 -4218
rect 2138 -4166 2190 -4156
rect 2138 -4228 2190 -4218
rect 1458 -4426 1622 -4390
rect 1662 -4276 1774 -4246
rect 1458 -4428 1510 -4426
rect 1458 -4490 1510 -4480
rect 1458 -4760 1494 -4490
rect 1578 -4520 1630 -4510
rect 1578 -4582 1630 -4572
rect 1460 -4802 1494 -4760
rect 1584 -4804 1620 -4582
rect 1662 -4672 1698 -4276
rect 2148 -4338 2182 -4228
rect 1740 -4376 2182 -4338
rect -396 -4876 1180 -4840
rect -396 -5084 -390 -4876
rect -396 -5120 1138 -5084
rect -396 -5456 -390 -5120
rect 1304 -5338 1340 -5068
rect 1382 -5234 1418 -5148
rect 1480 -5182 1698 -5148
rect 1374 -5244 1426 -5234
rect 1374 -5306 1426 -5296
rect 1296 -5348 1348 -5338
rect 1480 -5342 1514 -5182
rect 1654 -5244 1706 -5234
rect 1654 -5306 1706 -5296
rect 1296 -5410 1348 -5400
rect 1382 -5376 1514 -5342
rect -396 -5492 1138 -5456
rect -396 -5718 -390 -5492
rect 1382 -5494 1418 -5376
rect 1458 -5428 1510 -5418
rect 1458 -5490 1510 -5480
rect 1458 -5606 1494 -5490
rect 1662 -5492 1698 -5306
rect 1740 -5324 1776 -4376
rect 1804 -4428 1856 -4418
rect 1804 -4486 1856 -4480
rect 1804 -5296 1854 -4486
rect 3628 -4840 3634 -3652
rect 1918 -4876 3634 -4840
rect 3628 -5084 3634 -4876
rect 1942 -5120 3634 -5084
rect 1734 -5334 1786 -5324
rect 1734 -5396 1786 -5386
rect 1814 -5424 1854 -5296
rect -396 -5754 1176 -5718
rect -396 -6600 -390 -5754
rect 178 -6094 230 -6084
rect 1338 -6124 1374 -5952
rect 1584 -6028 1620 -5792
rect 1706 -6004 1742 -5792
rect 1804 -6004 1854 -5424
rect 3628 -5456 3634 -5120
rect 1942 -5492 3634 -5456
rect 3628 -5714 3634 -5492
rect 1910 -5750 3634 -5714
rect 1576 -6038 1628 -6028
rect 1706 -6040 1854 -6004
rect 1576 -6100 1628 -6090
rect 178 -6156 230 -6146
rect 1330 -6134 1382 -6124
rect 190 -6224 218 -6156
rect 1584 -6150 1620 -6100
rect 2576 -6134 2628 -6124
rect 1584 -6182 2342 -6150
rect 1330 -6196 1382 -6186
rect 150 -6252 2114 -6224
rect -396 -6636 54 -6600
rect -396 -6856 -390 -6636
rect -396 -6892 18 -6856
rect -396 -7228 -390 -6892
rect -396 -7264 18 -7228
rect -396 -7484 -390 -7264
rect -396 -7520 60 -7484
rect -396 -8105 -390 -7520
rect 150 -8016 178 -6252
rect 254 -6324 306 -6314
rect 254 -6386 306 -6376
rect 534 -6324 586 -6314
rect 534 -6386 586 -6376
rect 262 -6476 298 -6386
rect 542 -6476 578 -6386
rect 966 -6440 994 -6252
rect 1374 -6324 1426 -6314
rect 1374 -6386 1426 -6376
rect 1654 -6324 1706 -6314
rect 1654 -6386 1706 -6376
rect 822 -6476 1138 -6440
rect 1382 -6476 1418 -6386
rect 1662 -6476 1698 -6386
rect 2086 -6440 2114 -6252
rect 1942 -6476 2258 -6440
rect 212 -7020 246 -6900
rect 346 -6948 382 -6682
rect 338 -6958 390 -6948
rect 338 -7020 390 -7010
rect 212 -7030 298 -7020
rect 212 -7082 246 -7030
rect 212 -7092 298 -7082
rect 492 -7028 526 -6900
rect 626 -6948 662 -6682
rect 618 -6958 670 -6948
rect 618 -7020 670 -7010
rect 772 -7028 806 -6900
rect 492 -7038 544 -7028
rect 212 -7224 246 -7092
rect 492 -7100 544 -7090
rect 772 -7038 824 -7028
rect 772 -7100 824 -7090
rect 338 -7114 390 -7104
rect 338 -7176 390 -7166
rect 346 -7442 382 -7176
rect 492 -7224 526 -7100
rect 618 -7114 670 -7104
rect 618 -7176 670 -7166
rect 626 -7442 662 -7176
rect 772 -7224 806 -7100
rect 906 -7104 942 -6682
rect 1052 -7028 1086 -6900
rect 1052 -7038 1104 -7028
rect 1052 -7100 1104 -7090
rect 898 -7114 950 -7104
rect 898 -7176 950 -7166
rect 1052 -7224 1086 -7100
rect 1186 -7104 1222 -6682
rect 1332 -7028 1366 -6900
rect 1466 -6948 1502 -6682
rect 1458 -6958 1510 -6948
rect 1458 -7020 1510 -7010
rect 1612 -7028 1646 -6900
rect 1746 -6948 1782 -6682
rect 1738 -6958 1790 -6948
rect 1738 -7020 1790 -7010
rect 1892 -7028 1926 -6900
rect 1332 -7038 1384 -7028
rect 1332 -7100 1384 -7090
rect 1612 -7038 1664 -7028
rect 1612 -7100 1664 -7090
rect 1892 -7038 1944 -7028
rect 1892 -7100 1944 -7090
rect 1178 -7114 1230 -7104
rect 1178 -7176 1230 -7166
rect 1332 -7224 1366 -7100
rect 1458 -7114 1510 -7104
rect 1458 -7176 1510 -7166
rect 1466 -7442 1502 -7176
rect 1612 -7224 1646 -7100
rect 1738 -7114 1790 -7104
rect 1738 -7176 1790 -7166
rect 1746 -7442 1782 -7176
rect 1892 -7224 1926 -7100
rect 2026 -7104 2062 -6682
rect 2172 -7028 2206 -6900
rect 2172 -7038 2224 -7028
rect 2172 -7100 2224 -7090
rect 2018 -7114 2070 -7104
rect 2018 -7176 2070 -7166
rect 2172 -7224 2206 -7100
rect 2306 -7104 2342 -6182
rect 2576 -6196 2628 -6186
rect 2494 -6324 2546 -6314
rect 2494 -6386 2546 -6376
rect 2502 -6476 2538 -6386
rect 2586 -6732 2624 -6196
rect 2774 -6324 2826 -6314
rect 2774 -6386 2826 -6376
rect 2782 -6476 2818 -6386
rect 3628 -6408 3634 -5750
rect 3062 -6444 3634 -6408
rect 3628 -6662 3634 -6444
rect 2452 -7028 2486 -6900
rect 2586 -6948 2622 -6732
rect 2578 -6958 2630 -6948
rect 2578 -7020 2630 -7010
rect 2452 -7038 2504 -7028
rect 2732 -7048 2766 -6900
rect 2866 -6948 2902 -6682
rect 3030 -6698 3634 -6662
rect 2858 -6958 2910 -6948
rect 2858 -7020 2910 -7010
rect 3628 -7046 3634 -6698
rect 3478 -7048 3634 -7046
rect 2504 -7076 3634 -7048
rect 2452 -7100 2504 -7090
rect 2298 -7114 2350 -7104
rect 2298 -7176 2350 -7166
rect 2452 -7224 2486 -7100
rect 2578 -7114 2630 -7104
rect 2578 -7176 2630 -7166
rect 2586 -7442 2622 -7176
rect 2732 -7224 2766 -7076
rect 2858 -7114 2910 -7104
rect 2858 -7176 2910 -7166
rect 2866 -7442 2902 -7176
rect 3628 -7358 3634 -7076
rect 3032 -7394 3634 -7358
rect 262 -7684 578 -7648
rect 406 -8016 434 -7684
rect 822 -7738 858 -7684
rect 814 -7748 866 -7738
rect 814 -7810 866 -7800
rect 906 -7832 942 -7442
rect 1102 -7738 1138 -7684
rect 1094 -7748 1146 -7738
rect 1094 -7810 1146 -7800
rect 1186 -7832 1222 -7442
rect 1382 -7684 1698 -7648
rect 898 -7842 950 -7832
rect 898 -7904 950 -7894
rect 1178 -7842 1230 -7832
rect 1178 -7904 1230 -7894
rect 1526 -8016 1554 -7684
rect 1942 -7738 1978 -7684
rect 1934 -7748 1986 -7738
rect 1934 -7810 1986 -7800
rect 2026 -7832 2062 -7442
rect 2222 -7738 2258 -7684
rect 2214 -7748 2266 -7738
rect 2214 -7810 2266 -7800
rect 2306 -7832 2342 -7442
rect 3628 -7616 3634 -7394
rect 2502 -7684 2818 -7648
rect 3062 -7652 3634 -7616
rect 2018 -7842 2070 -7832
rect 2018 -7904 2070 -7894
rect 2298 -7842 2350 -7832
rect 2298 -7904 2350 -7894
rect 2646 -8016 2674 -7684
rect 150 -8044 2674 -8016
rect -502 -8416 -390 -8105
rect 3628 -8105 3634 -7652
rect 3734 -8105 3740 -2395
rect 210 -8416 220 -8116
rect 3018 -8416 3028 -8116
rect 3628 -8416 3740 -8105
rect -502 -8422 3740 -8416
rect -502 -8522 -396 -8422
rect 3634 -8522 3740 -8422
rect -502 -8528 3740 -8522
<< via1 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -110 440 -58 492
rect 170 440 222 492
rect -26 346 26 398
rect 60 -382 112 -330
rect -26 -1114 26 -1062
rect 450 440 502 492
rect 254 346 306 398
rect 340 -382 392 -330
rect 730 440 782 492
rect 534 346 586 398
rect 620 -382 672 -330
rect 1010 440 1062 492
rect 814 346 866 398
rect 900 -382 952 -330
rect 1290 440 1342 492
rect 1094 346 1146 398
rect 1180 -382 1232 -330
rect 1570 440 1622 492
rect 1374 346 1426 398
rect 1460 -382 1512 -330
rect 1850 440 1902 492
rect 1654 346 1706 398
rect 1740 -382 1792 -330
rect 2130 440 2182 492
rect 1934 346 1986 398
rect 2020 -382 2072 -330
rect 2410 440 2462 492
rect 2214 346 2266 398
rect 2300 -382 2352 -330
rect 2690 440 2742 492
rect 2494 346 2546 398
rect 2580 -382 2632 -330
rect 2970 440 3022 492
rect 2774 346 2826 398
rect 2860 -382 2912 -330
rect 3238 238 3290 290
rect 3520 238 3572 290
rect 3140 -382 3192 -330
rect 254 -1114 306 -1062
rect 534 -1114 586 -1062
rect 814 -1114 866 -1062
rect 1094 -1114 1146 -1062
rect 1934 -1114 1986 -1062
rect 2214 -1114 2266 -1062
rect 2494 -1114 2546 -1062
rect 2774 -1114 2826 -1062
rect 3054 -1114 3106 -1062
rect 1374 -1230 1426 -1178
rect 1654 -1230 1706 -1178
rect 414 -1514 466 -1462
rect 2478 -1424 2530 -1372
rect 900 -2194 952 -2142
rect 2774 -2186 2826 -2134
rect 330 -2274 382 -2222
rect 610 -2274 662 -2222
rect 178 -2374 230 -2322
rect 254 -2474 306 -2422
rect 458 -2374 510 -2322
rect 534 -2474 586 -2422
rect 814 -2474 866 -2422
rect 1450 -2274 1502 -2222
rect 1730 -2274 1782 -2222
rect 2570 -2274 2622 -2222
rect 1298 -2374 1350 -2322
rect 1094 -2474 1146 -2422
rect 1374 -2474 1426 -2422
rect 1578 -2374 1630 -2322
rect 1654 -2474 1706 -2422
rect 2418 -2374 2470 -2322
rect 1934 -2474 1986 -2422
rect 2214 -2474 2266 -2422
rect 2494 -2474 2546 -2422
rect 2698 -2374 2750 -2322
rect 2850 -2274 2902 -2222
rect 2774 -2474 2826 -2422
rect 178 -3198 230 -3146
rect 458 -3198 510 -3146
rect 738 -3194 790 -3142
rect 330 -3298 382 -3246
rect 1018 -3194 1070 -3142
rect 1298 -3198 1350 -3146
rect 1578 -3198 1630 -3146
rect 1858 -3194 1910 -3142
rect 610 -3298 662 -3246
rect 890 -3298 942 -3246
rect 1170 -3298 1222 -3246
rect 1450 -3298 1502 -3246
rect 254 -4018 306 -3966
rect 534 -4018 586 -3966
rect 814 -4018 866 -3966
rect 890 -4118 942 -4066
rect 1094 -4018 1146 -3966
rect 1374 -4018 1426 -3966
rect 1170 -4118 1222 -4066
rect 738 -4218 790 -4166
rect 1018 -4218 1070 -4166
rect 2138 -3194 2190 -3142
rect 2418 -3198 2470 -3146
rect 2698 -3198 2750 -3146
rect 1730 -3298 1782 -3246
rect 2010 -3298 2062 -3246
rect 2290 -3298 2342 -3246
rect 2570 -3298 2622 -3246
rect 2850 -3298 2902 -3246
rect 1654 -4018 1706 -3966
rect 1934 -4018 1986 -3966
rect 2010 -4118 2062 -4066
rect 2214 -4018 2266 -3966
rect 2494 -4018 2546 -3966
rect 2774 -4018 2826 -3966
rect 2290 -4118 2342 -4066
rect 1858 -4218 1910 -4166
rect 2138 -4218 2190 -4166
rect 1458 -4480 1510 -4428
rect 1578 -4572 1630 -4520
rect 1374 -5296 1426 -5244
rect 1654 -5296 1706 -5244
rect 1296 -5400 1348 -5348
rect 1458 -5480 1510 -5428
rect 1804 -4480 1856 -4428
rect 1734 -5386 1786 -5334
rect 178 -6146 230 -6094
rect 1576 -6090 1628 -6038
rect 1330 -6186 1382 -6134
rect 254 -6376 306 -6324
rect 534 -6376 586 -6324
rect 1374 -6376 1426 -6324
rect 1654 -6376 1706 -6324
rect 338 -7010 390 -6958
rect 246 -7082 298 -7030
rect 618 -7010 670 -6958
rect 492 -7090 544 -7038
rect 772 -7090 824 -7038
rect 338 -7166 390 -7114
rect 618 -7166 670 -7114
rect 1052 -7090 1104 -7038
rect 898 -7166 950 -7114
rect 1458 -7010 1510 -6958
rect 1738 -7010 1790 -6958
rect 1332 -7090 1384 -7038
rect 1612 -7090 1664 -7038
rect 1892 -7090 1944 -7038
rect 1178 -7166 1230 -7114
rect 1458 -7166 1510 -7114
rect 1738 -7166 1790 -7114
rect 2172 -7090 2224 -7038
rect 2018 -7166 2070 -7114
rect 2576 -6186 2628 -6134
rect 2494 -6376 2546 -6324
rect 2774 -6376 2826 -6324
rect 2578 -7010 2630 -6958
rect 2452 -7090 2504 -7038
rect 2858 -7010 2910 -6958
rect 2298 -7166 2350 -7114
rect 2578 -7166 2630 -7114
rect 2858 -7166 2910 -7114
rect 814 -7800 866 -7748
rect 1094 -7800 1146 -7748
rect 898 -7894 950 -7842
rect 1178 -7894 1230 -7842
rect 1934 -7800 1986 -7748
rect 2214 -7800 2266 -7748
rect 2018 -7894 2070 -7842
rect 2298 -7894 2350 -7842
rect -390 -8416 210 -8116
rect 3028 -8416 3628 -8116
<< metal2 >>
rect -390 1016 210 1026
rect -390 706 210 716
rect 3028 1016 3628 1026
rect 3028 706 3628 716
rect -120 440 -110 492
rect -58 440 170 492
rect 222 440 450 492
rect 502 440 730 492
rect 782 440 1010 492
rect 1062 440 1290 492
rect 1342 440 1570 492
rect 1622 440 1850 492
rect 1902 440 2130 492
rect 2182 440 2410 492
rect 2462 440 2690 492
rect 2742 440 2970 492
rect 3022 440 3032 492
rect -290 346 -26 398
rect 26 346 36 398
rect 244 346 254 398
rect 306 396 316 398
rect 524 396 534 398
rect 306 346 534 396
rect 586 396 596 398
rect 804 396 814 398
rect 586 346 814 396
rect 866 396 876 398
rect 1084 396 1094 398
rect 866 346 1094 396
rect 1146 396 1156 398
rect 1364 396 1374 398
rect 1146 346 1374 396
rect 1426 396 1436 398
rect 1644 396 1654 398
rect 1426 346 1654 396
rect 1706 396 1716 398
rect 1924 396 1934 398
rect 1706 346 1934 396
rect 1986 396 1996 398
rect 2204 396 2214 398
rect 1986 346 2214 396
rect 2266 396 2276 398
rect 2484 396 2494 398
rect 2266 346 2494 396
rect 2546 396 2556 398
rect 2764 396 2774 398
rect 2546 346 2774 396
rect 2826 396 2836 398
rect 3338 396 3390 398
rect 2826 346 3390 396
rect -290 298 -138 346
rect -190 -1178 -138 298
rect 3238 290 3290 300
rect 50 -382 60 -330
rect 112 -382 340 -330
rect 392 -382 620 -330
rect 672 -382 900 -330
rect 952 -382 1180 -330
rect 1232 -382 1460 -330
rect 1512 -382 1522 -330
rect 1730 -382 1740 -330
rect 1792 -382 2020 -330
rect 2072 -382 2300 -330
rect 2352 -382 2580 -330
rect 2632 -382 2860 -330
rect 2912 -382 3140 -330
rect 3192 -382 3202 -330
rect -36 -1114 -26 -1062
rect 26 -1114 254 -1062
rect 306 -1114 534 -1062
rect 586 -1114 814 -1062
rect 866 -1114 1094 -1062
rect 1146 -1114 1934 -1062
rect 1986 -1114 2214 -1062
rect 2266 -1114 2494 -1062
rect 2546 -1114 2774 -1062
rect 2826 -1114 3054 -1062
rect 3106 -1114 3116 -1062
rect -190 -1230 1374 -1178
rect 1426 -1230 1436 -1178
rect 414 -1462 466 -1452
rect 414 -1764 466 -1514
rect 964 -1466 1016 -1230
rect 1514 -1258 1566 -1114
rect 3238 -1178 3290 238
rect 1644 -1230 1654 -1178
rect 1706 -1230 3290 -1178
rect 3338 -1258 3390 346
rect 3498 300 3598 400
rect 3520 290 3572 300
rect 3520 232 3572 238
rect 1514 -1310 3390 -1258
rect 2478 -1372 2530 -1362
rect 1954 -1466 2000 -1464
rect 2478 -1466 2530 -1424
rect 964 -1518 2530 -1466
rect 414 -1804 806 -1764
rect 774 -2154 806 -1804
rect 890 -2154 900 -2142
rect 774 -2194 900 -2154
rect 952 -2194 962 -2142
rect 1954 -2222 2000 -1518
rect 2916 -1792 2972 -1310
rect 2894 -1892 2994 -1792
rect 2916 -2134 2972 -1892
rect 2764 -2186 2774 -2134
rect 2826 -2186 2972 -2134
rect 2916 -2188 2972 -2186
rect 320 -2274 330 -2222
rect 382 -2274 610 -2222
rect 662 -2274 1450 -2222
rect 1502 -2274 1730 -2222
rect 1782 -2274 2570 -2222
rect 2622 -2274 2850 -2222
rect 2902 -2274 3104 -2222
rect -76 -2374 178 -2322
rect 230 -2374 458 -2322
rect 510 -2374 1298 -2322
rect 1350 -2374 1578 -2322
rect 1630 -2374 2418 -2322
rect 2470 -2374 2698 -2322
rect 2750 -2374 2760 -2322
rect -76 -4166 -24 -2374
rect 58 -2474 254 -2422
rect 306 -2474 534 -2422
rect 586 -2474 814 -2422
rect 866 -2474 1094 -2422
rect 1146 -2474 1374 -2422
rect 1426 -2474 1654 -2422
rect 1706 -2474 1934 -2422
rect 1986 -2474 2214 -2422
rect 2266 -2474 2494 -2422
rect 2546 -2474 2774 -2422
rect 2826 -2474 3022 -2422
rect 58 -3966 110 -2474
rect 728 -3146 738 -3142
rect 168 -3198 178 -3146
rect 230 -3198 458 -3146
rect 510 -3194 738 -3146
rect 790 -3146 800 -3142
rect 1008 -3146 1018 -3142
rect 790 -3194 1018 -3146
rect 1070 -3146 1080 -3142
rect 1848 -3146 1858 -3142
rect 1070 -3194 1298 -3146
rect 510 -3198 1298 -3194
rect 1350 -3198 1578 -3146
rect 1630 -3194 1858 -3146
rect 1910 -3146 1920 -3142
rect 2128 -3146 2138 -3142
rect 1910 -3194 2138 -3146
rect 2190 -3146 2200 -3142
rect 2190 -3194 2418 -3146
rect 1630 -3198 2418 -3194
rect 2470 -3198 2698 -3146
rect 2750 -3198 2760 -3146
rect 320 -3298 330 -3246
rect 382 -3298 610 -3246
rect 662 -3298 890 -3246
rect 942 -3298 1170 -3246
rect 1222 -3298 1450 -3246
rect 1502 -3298 1730 -3246
rect 1782 -3298 2010 -3246
rect 2062 -3298 2290 -3246
rect 2342 -3298 2570 -3246
rect 2622 -3298 2850 -3246
rect 2902 -3298 2912 -3246
rect 330 -3300 2902 -3298
rect 2970 -3966 3022 -2474
rect 58 -4018 254 -3966
rect 306 -4018 534 -3966
rect 586 -4018 814 -3966
rect 866 -4018 1094 -3966
rect 1146 -4018 1374 -3966
rect 1426 -4018 1654 -3966
rect 1706 -4018 1934 -3966
rect 1986 -4018 2214 -3966
rect 2266 -4018 2494 -3966
rect 2546 -4018 2774 -3966
rect 2826 -4018 3022 -3966
rect 3052 -4066 3104 -2274
rect 880 -4118 890 -4066
rect 942 -4118 1170 -4066
rect 1222 -4118 2010 -4066
rect 2062 -4118 2290 -4066
rect 2342 -4118 3104 -4066
rect -76 -4218 738 -4166
rect 790 -4218 1018 -4166
rect 1070 -4218 1858 -4166
rect 1910 -4218 2138 -4166
rect 2190 -4218 2200 -4166
rect 1448 -4480 1458 -4428
rect 1510 -4480 1804 -4428
rect 1856 -4480 1866 -4428
rect 1568 -4572 1578 -4520
rect 1630 -4572 1876 -4520
rect 1364 -5296 1374 -5244
rect 1426 -5296 1654 -5244
rect 1706 -5296 1716 -5244
rect 1724 -5346 1734 -5334
rect 1286 -5400 1296 -5348
rect 1348 -5400 1358 -5348
rect 1554 -5380 1734 -5346
rect 1296 -6038 1348 -5400
rect 1554 -5428 1588 -5380
rect 1724 -5386 1734 -5380
rect 1786 -5386 1796 -5334
rect 1448 -5480 1458 -5428
rect 1510 -5480 1588 -5428
rect -152 -6094 -52 -6060
rect 1296 -6090 1576 -6038
rect 1628 -6090 1638 -6038
rect -152 -6146 178 -6094
rect 230 -6146 240 -6094
rect 1826 -6134 1876 -4572
rect -152 -6160 -52 -6146
rect 1320 -6186 1330 -6134
rect 1382 -6186 2576 -6134
rect 2628 -6186 2638 -6134
rect 2836 -6324 2936 -6276
rect 138 -6376 254 -6324
rect 306 -6376 534 -6324
rect 586 -6376 1374 -6324
rect 1426 -6376 1654 -6324
rect 1706 -6376 2494 -6324
rect 2546 -6376 2774 -6324
rect 2826 -6376 2936 -6324
rect 138 -7748 196 -6376
rect 328 -7010 338 -6958
rect 390 -7010 618 -6958
rect 670 -7010 1458 -6958
rect 1510 -7010 1738 -6958
rect 1790 -7010 2578 -6958
rect 2630 -7010 2858 -6958
rect 2910 -7010 3026 -6958
rect 236 -7082 246 -7030
rect 298 -7048 308 -7030
rect 482 -7048 492 -7038
rect 298 -7076 492 -7048
rect 298 -7082 308 -7076
rect 482 -7090 492 -7076
rect 544 -7048 554 -7038
rect 762 -7048 772 -7038
rect 544 -7076 772 -7048
rect 544 -7090 554 -7076
rect 762 -7090 772 -7076
rect 824 -7048 834 -7038
rect 1042 -7048 1052 -7038
rect 824 -7076 1052 -7048
rect 824 -7090 834 -7076
rect 1042 -7090 1052 -7076
rect 1104 -7048 1114 -7038
rect 1322 -7048 1332 -7038
rect 1104 -7076 1332 -7048
rect 1104 -7090 1114 -7076
rect 1322 -7090 1332 -7076
rect 1384 -7048 1394 -7038
rect 1602 -7048 1612 -7038
rect 1384 -7076 1612 -7048
rect 1384 -7090 1394 -7076
rect 1602 -7090 1612 -7076
rect 1664 -7048 1674 -7038
rect 1882 -7048 1892 -7038
rect 1664 -7076 1892 -7048
rect 1664 -7090 1674 -7076
rect 1882 -7090 1892 -7076
rect 1944 -7048 1954 -7038
rect 2162 -7048 2172 -7038
rect 1944 -7076 2172 -7048
rect 1944 -7090 1954 -7076
rect 2162 -7090 2172 -7076
rect 2224 -7048 2234 -7038
rect 2442 -7048 2452 -7038
rect 2224 -7076 2452 -7048
rect 2224 -7090 2234 -7076
rect 2442 -7090 2452 -7076
rect 2504 -7090 2514 -7038
rect 328 -7166 338 -7114
rect 390 -7118 396 -7114
rect 612 -7118 618 -7114
rect 390 -7166 618 -7118
rect 670 -7118 676 -7114
rect 892 -7118 898 -7114
rect 670 -7166 898 -7118
rect 950 -7118 956 -7114
rect 1172 -7118 1178 -7114
rect 950 -7166 1178 -7118
rect 1230 -7118 1236 -7114
rect 1452 -7118 1458 -7114
rect 1230 -7166 1458 -7118
rect 1510 -7118 1516 -7114
rect 1732 -7118 1738 -7114
rect 1510 -7166 1738 -7118
rect 1790 -7118 1796 -7114
rect 2012 -7118 2018 -7114
rect 1790 -7166 2018 -7118
rect 2070 -7118 2076 -7114
rect 2292 -7118 2298 -7114
rect 2070 -7166 2298 -7118
rect 2350 -7118 2356 -7114
rect 2572 -7118 2578 -7114
rect 2350 -7166 2578 -7118
rect 2630 -7118 2636 -7114
rect 2852 -7118 2858 -7114
rect 2630 -7166 2858 -7118
rect 2910 -7166 2920 -7114
rect 138 -7800 814 -7748
rect 866 -7800 1094 -7748
rect 1146 -7800 1934 -7748
rect 1986 -7800 2214 -7748
rect 2266 -7800 2276 -7748
rect 2978 -7842 3026 -7010
rect 888 -7894 898 -7842
rect 950 -7894 1178 -7842
rect 1230 -7894 2018 -7842
rect 2070 -7894 2298 -7842
rect 2350 -7894 3026 -7842
rect -390 -8116 210 -8106
rect -390 -8426 210 -8416
rect 3028 -8116 3628 -8106
rect 3028 -8426 3628 -8416
<< via2 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -390 -8416 210 -8116
rect 3028 -8416 3628 -8116
<< metal3 >>
rect -400 1016 220 1021
rect -400 716 -390 1016
rect 210 716 220 1016
rect -400 711 220 716
rect 3018 1016 3638 1021
rect 3018 716 3028 1016
rect 3628 716 3638 1016
rect 3018 711 3638 716
rect -400 -8116 220 -8111
rect -400 -8416 -390 -8116
rect 210 -8416 220 -8116
rect -400 -8421 220 -8416
rect 3018 -8116 3638 -8111
rect 3018 -8416 3028 -8116
rect 3628 -8416 3638 -8116
rect 3018 -8421 3638 -8416
<< via3 >>
rect -390 716 210 1016
rect 3028 716 3628 1016
rect -390 -8416 210 -8116
rect 3028 -8416 3628 -8116
<< metal4 >>
rect -391 1016 211 1017
rect -391 716 -390 1016
rect 210 716 211 1016
rect -391 715 211 716
rect 3027 1016 3629 1017
rect 3027 716 3028 1016
rect 3628 716 3629 1016
rect 3027 715 3629 716
rect -391 -8116 211 -8115
rect -391 -8416 -390 -8116
rect 210 -8416 211 -8116
rect -391 -8417 211 -8416
rect 3027 -8116 3629 -8115
rect 3027 -8416 3028 -8116
rect 3628 -8416 3629 -8116
rect 3027 -8417 3629 -8416
use sky130_fd_pr__nfet_01v8_7B6TAC  sky130_fd_pr__nfet_01v8_7B6TAC_0 
timestamp 1733619730
transform 1 0 3080 0 1 -7410
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PHZV97  sky130_fd_pr__nfet_01v8_PHZV97_0 
timestamp 1733217049
transform 1 0 1399 0 1 -4909
box -99 -288 99 288
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm1 
timestamp 1733217602
transform 1 0 0 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm2
timestamp 1733217602
transform 1 0 280 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm3
timestamp 1733217602
transform 1 0 560 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm4
timestamp 1733217602
transform 1 0 840 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm5
timestamp 1733217602
transform 1 0 1120 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm6
timestamp 1733217602
transform 1 0 1400 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm7
timestamp 1733217602
transform 1 0 1680 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm8
timestamp 1733217602
transform 1 0 1960 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm9
timestamp 1733217602
transform 1 0 2240 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm10
timestamp 1733217602
transform 1 0 2520 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm11
timestamp 1733217602
transform 1 0 2800 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm12
timestamp 1733217602
transform 1 0 3080 0 1 0
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm13
timestamp 1733217602
transform 1 0 0 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm14
timestamp 1733217602
transform 1 0 280 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm15
timestamp 1733217602
transform 1 0 560 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm16
timestamp 1733217602
transform 1 0 840 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm17
timestamp 1733217602
transform 1 0 1120 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm18
timestamp 1733217602
transform 1 0 1400 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm19
timestamp 1733217602
transform 1 0 1680 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm20
timestamp 1733217602
transform 1 0 1960 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm21
timestamp 1733217602
transform 1 0 2240 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm22
timestamp 1733217602
transform 1 0 2520 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm23
timestamp 1733217602
transform 1 0 2800 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__pfet_01v8_MJ75SZ  xm24
timestamp 1733217602
transform 1 0 3080 0 1 -716
box -109 -300 109 300
use sky130_fd_pr__nfet_01v8_PHZV97  xm25
timestamp 1733217049
transform 1 0 279 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm26
timestamp 1733217049
transform 1 0 559 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm27
timestamp 1733217049
transform 1 0 839 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm28
timestamp 1733217049
transform 1 0 1119 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm29
timestamp 1733217049
transform 1 0 1399 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm30
timestamp 1733217049
transform 1 0 1679 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm31
timestamp 1733217049
transform 1 0 1959 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm32
timestamp 1733217049
transform 1 0 2239 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm33
timestamp 1733217049
transform 1 0 2519 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm34
timestamp 1733217049
transform 1 0 2799 0 1 -2809
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm35
timestamp 1733217049
transform 1 0 279 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm36
timestamp 1733217049
transform 1 0 559 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm37
timestamp 1733217049
transform 1 0 839 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm38
timestamp 1733217049
transform 1 0 1119 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm39
timestamp 1733217049
transform 1 0 1399 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm40
timestamp 1733217049
transform 1 0 1679 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm41
timestamp 1733217049
transform 1 0 1959 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm42
timestamp 1733217049
transform 1 0 2239 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm43
timestamp 1733217049
transform 1 0 2519 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm44
timestamp 1733217049
transform 1 0 2799 0 1 -3629
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_PHZV97  xm46
timestamp 1733217049
transform 1 0 1679 0 1 -4909
box -99 -288 99 288
use sky130_fd_pr__nfet_01v8_72KZQ8  xm47 
timestamp 1733216309
transform 1 0 1398 0 1 -5736
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm48
timestamp 1733216309
transform 1 0 1678 0 1 -5736
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm49
timestamp 1733216309
transform 1 0 279 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm50
timestamp 1733216309
transform 1 0 559 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm51
timestamp 1733216309
transform 1 0 839 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm52
timestamp 1733216309
transform 1 0 1119 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm53
timestamp 1733216309
transform 1 0 1399 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm54
timestamp 1733216309
transform 1 0 1679 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm55
timestamp 1733216309
transform 1 0 1959 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm56
timestamp 1733216309
transform 1 0 2239 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm57
timestamp 1733216309
transform 1 0 2519 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm58
timestamp 1733216309
transform 1 0 2799 0 1 -6681
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm59 
timestamp 1733216309
transform 1 0 279 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm60
timestamp 1733216309
transform 1 0 559 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm61
timestamp 1733216309
transform 1 0 839 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm62
timestamp 1733216309
transform 1 0 1119 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm63
timestamp 1733216309
transform 1 0 1399 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm64
timestamp 1733216309
transform 1 0 1679 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm65
timestamp 1733216309
transform 1 0 1959 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm66
timestamp 1733216309
transform 1 0 2239 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm67
timestamp 1733216309
transform 1 0 2519 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm68
timestamp 1733216309
transform 1 0 2799 0 1 -7441
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm69
timestamp 1733216309
transform 1 0 0 0 1 -2778
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm70
timestamp 1733216309
transform 1 0 0 0 1 -3598
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm71
timestamp 1733216309
transform 1 0 3080 0 1 -2778
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm72
timestamp 1733216309
transform 1 0 3080 0 1 -3598
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm73
timestamp 1733216309
transform 1 0 0 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm74
timestamp 1733216309
transform 1 0 0 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm75
timestamp 1733216309
transform 1 0 280 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm76
timestamp 1733216309
transform 1 0 280 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm77
timestamp 1733216309
transform 1 0 560 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm78
timestamp 1733216309
transform 1 0 560 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm79
timestamp 1733216309
transform 1 0 840 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm80
timestamp 1733216309
transform 1 0 840 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm81
timestamp 1733216309
transform 1 0 1120 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm82
timestamp 1733216309
transform 1 0 1120 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm83
timestamp 1733216309
transform 1 0 1960 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm84
timestamp 1733216309
transform 1 0 1960 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm85
timestamp 1733216309
transform 1 0 2240 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm86
timestamp 1733216309
transform 1 0 2240 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm87
timestamp 1733216309
transform 1 0 2520 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm88
timestamp 1733216309
transform 1 0 2520 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm89
timestamp 1733216309
transform 1 0 2800 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm90
timestamp 1733216309
transform 1 0 2800 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm91
timestamp 1733216309
transform 1 0 3080 0 1 -4878
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm92
timestamp 1733216309
transform 1 0 3080 0 1 -5698
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_PRFKA7  xm93
timestamp 1733216309
transform 1 0 0 0 1 -6650
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm94
timestamp 1733216309
transform 1 0 0 0 1 -7470
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_72KZQ8  xm95
timestamp 1733216309
transform 1 0 3080 0 1 -6650
box -73 -257 73 257
<< labels >>
rlabel via1 -146 874 -46 974 1 VDD
port 1 n
rlabel metal2 -290 298 -190 398 1 Voutminus
port 9 n
rlabel metal2 3498 300 3598 400 1 Voutplus
port 10 n
rlabel metal2 2894 -1892 2994 -1792 1 CLK
port 11 n
rlabel via1 3262 -8306 3362 -8206 1 VSS
port 8 n
rlabel metal2 -152 -6160 -52 -6060 1 Vioplus
port 12 n
rlabel metal2 2836 -6376 2936 -6276 1 Viominus
port 13 n
<< properties >>
string FIXED_BBOX -446 -8472 3684 -2028
<< end >>
