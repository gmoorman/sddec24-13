* NGSPICE file created from 2x2.ext - technology: sky130B

.subckt sky130_fd_pr_reram__reram_cell_X TE BE
X0 TE BE sky130_fd_pr_reram__reram_cell area_ox=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B a_50_n700# a_n242_n922# a_n108_n700# a_n50_n788#
X0 a_50_n700# a_n50_n788# a_n108_n700# a_n242_n922# sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=0.5
.ends

.subckt x1T1R SL WL BL VSS
XXR1 BL XR1/BE sky130_fd_pr_reram__reram_cell_X
XXM1 XR1/BE VSS SL WL sky130_fd_pr__nfet_g5v0d10v5_9YEQ2B
.ends

.subckt x2x2 BL2 BL1 VSS WL1 WL2 SL1 SL2
Xx1 SL1 WL1 BL1 VSS x1T1R
Xx3 SL2 WL2 BL1 VSS x1T1R
Xx2 SL1 WL1 BL2 VSS x1T1R
Xx4 SL2 WL2 BL2 VSS x1T1R
.ends

